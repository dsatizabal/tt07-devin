VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_devin
  CLASS BLOCK ;
  FOREIGN tt_um_devin ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.300000 ;
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER met4 ;
        RECT 156.410 0.000 157.310 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.300000 ;
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER met4 ;
        RECT 134.330 0.000 135.230 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.250 0.000 113.150 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.170 0.000 91.070 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.090 0.000 68.990 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.010 0.000 46.910 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.930 0.000 24.830 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1.850 0.000 2.750 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 340.199982 ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 131.500 1.750 134.600 211.700 ;
      LAYER nwell ;
        RECT 134.800 1.760 137.990 211.710 ;
      LAYER pwell ;
        RECT 153.550 1.760 156.650 211.770 ;
      LAYER nwell ;
        RECT 156.850 1.770 160.040 211.780 ;
      LAYER li1 ;
        RECT 131.680 211.450 134.420 211.520 ;
        RECT 131.550 211.350 134.420 211.450 ;
        RECT 131.550 209.940 131.850 211.350 ;
        RECT 132.190 210.480 132.360 210.810 ;
        RECT 132.530 210.780 133.570 210.950 ;
        RECT 132.530 210.340 133.570 210.510 ;
        RECT 133.740 210.480 133.910 210.810 ;
        RECT 134.250 209.940 134.420 211.350 ;
        RECT 131.550 209.800 134.420 209.940 ;
        RECT 131.680 209.770 134.420 209.800 ;
        RECT 134.980 211.480 137.810 211.530 ;
        RECT 153.730 211.520 156.470 211.590 ;
        RECT 134.980 211.360 137.930 211.480 ;
        RECT 134.980 209.950 135.150 211.360 ;
        RECT 135.490 210.490 135.660 210.820 ;
        RECT 135.875 210.790 136.915 210.960 ;
        RECT 135.875 210.350 136.915 210.520 ;
        RECT 137.130 210.490 137.300 210.820 ;
        RECT 137.640 209.950 137.930 211.360 ;
        RECT 134.980 209.830 137.930 209.950 ;
        RECT 153.600 211.420 156.470 211.520 ;
        RECT 153.600 210.010 153.900 211.420 ;
        RECT 154.240 210.550 154.410 210.880 ;
        RECT 154.580 210.850 155.620 211.020 ;
        RECT 154.580 210.410 155.620 210.580 ;
        RECT 155.790 210.550 155.960 210.880 ;
        RECT 156.300 210.010 156.470 211.420 ;
        RECT 153.600 209.870 156.470 210.010 ;
        RECT 153.730 209.840 156.470 209.870 ;
        RECT 157.030 211.550 159.860 211.600 ;
        RECT 157.030 211.430 159.980 211.550 ;
        RECT 157.030 210.020 157.200 211.430 ;
        RECT 157.540 210.560 157.710 210.890 ;
        RECT 157.925 210.860 158.965 211.030 ;
        RECT 157.925 210.420 158.965 210.590 ;
        RECT 159.180 210.560 159.350 210.890 ;
        RECT 159.690 210.020 159.980 211.430 ;
        RECT 157.030 209.900 159.980 210.020 ;
        RECT 157.030 209.850 159.860 209.900 ;
        RECT 134.980 209.780 137.810 209.830 ;
        RECT 131.680 209.350 134.420 209.420 ;
        RECT 131.550 209.250 134.420 209.350 ;
        RECT 131.550 207.840 131.850 209.250 ;
        RECT 132.190 208.380 132.360 208.710 ;
        RECT 132.530 208.680 133.570 208.850 ;
        RECT 132.530 208.240 133.570 208.410 ;
        RECT 133.740 208.380 133.910 208.710 ;
        RECT 134.250 207.840 134.420 209.250 ;
        RECT 131.550 207.700 134.420 207.840 ;
        RECT 131.680 207.670 134.420 207.700 ;
        RECT 134.980 209.380 137.810 209.430 ;
        RECT 153.730 209.420 156.470 209.490 ;
        RECT 134.980 209.260 137.930 209.380 ;
        RECT 134.980 207.850 135.150 209.260 ;
        RECT 135.490 208.390 135.660 208.720 ;
        RECT 135.875 208.690 136.915 208.860 ;
        RECT 135.875 208.250 136.915 208.420 ;
        RECT 137.130 208.390 137.300 208.720 ;
        RECT 137.640 207.850 137.930 209.260 ;
        RECT 134.980 207.730 137.930 207.850 ;
        RECT 153.600 209.320 156.470 209.420 ;
        RECT 153.600 207.910 153.900 209.320 ;
        RECT 154.240 208.450 154.410 208.780 ;
        RECT 154.580 208.750 155.620 208.920 ;
        RECT 154.580 208.310 155.620 208.480 ;
        RECT 155.790 208.450 155.960 208.780 ;
        RECT 156.300 207.910 156.470 209.320 ;
        RECT 153.600 207.770 156.470 207.910 ;
        RECT 153.730 207.740 156.470 207.770 ;
        RECT 157.030 209.450 159.860 209.500 ;
        RECT 157.030 209.330 159.980 209.450 ;
        RECT 157.030 207.920 157.200 209.330 ;
        RECT 157.540 208.460 157.710 208.790 ;
        RECT 157.925 208.760 158.965 208.930 ;
        RECT 157.925 208.320 158.965 208.490 ;
        RECT 159.180 208.460 159.350 208.790 ;
        RECT 159.690 207.920 159.980 209.330 ;
        RECT 157.030 207.800 159.980 207.920 ;
        RECT 157.030 207.750 159.860 207.800 ;
        RECT 134.980 207.680 137.810 207.730 ;
        RECT 131.680 207.250 134.420 207.320 ;
        RECT 131.550 207.150 134.420 207.250 ;
        RECT 131.550 205.740 131.850 207.150 ;
        RECT 132.190 206.280 132.360 206.610 ;
        RECT 132.530 206.580 133.570 206.750 ;
        RECT 132.530 206.140 133.570 206.310 ;
        RECT 133.740 206.280 133.910 206.610 ;
        RECT 134.250 205.740 134.420 207.150 ;
        RECT 131.550 205.600 134.420 205.740 ;
        RECT 131.680 205.570 134.420 205.600 ;
        RECT 134.980 207.280 137.810 207.330 ;
        RECT 153.730 207.320 156.470 207.390 ;
        RECT 134.980 207.160 137.930 207.280 ;
        RECT 134.980 205.750 135.150 207.160 ;
        RECT 135.490 206.290 135.660 206.620 ;
        RECT 135.875 206.590 136.915 206.760 ;
        RECT 135.875 206.150 136.915 206.320 ;
        RECT 137.130 206.290 137.300 206.620 ;
        RECT 137.640 205.750 137.930 207.160 ;
        RECT 134.980 205.630 137.930 205.750 ;
        RECT 153.600 207.220 156.470 207.320 ;
        RECT 153.600 205.810 153.900 207.220 ;
        RECT 154.240 206.350 154.410 206.680 ;
        RECT 154.580 206.650 155.620 206.820 ;
        RECT 154.580 206.210 155.620 206.380 ;
        RECT 155.790 206.350 155.960 206.680 ;
        RECT 156.300 205.810 156.470 207.220 ;
        RECT 153.600 205.670 156.470 205.810 ;
        RECT 153.730 205.640 156.470 205.670 ;
        RECT 157.030 207.350 159.860 207.400 ;
        RECT 157.030 207.230 159.980 207.350 ;
        RECT 157.030 205.820 157.200 207.230 ;
        RECT 157.540 206.360 157.710 206.690 ;
        RECT 157.925 206.660 158.965 206.830 ;
        RECT 157.925 206.220 158.965 206.390 ;
        RECT 159.180 206.360 159.350 206.690 ;
        RECT 159.690 205.820 159.980 207.230 ;
        RECT 157.030 205.700 159.980 205.820 ;
        RECT 157.030 205.650 159.860 205.700 ;
        RECT 134.980 205.580 137.810 205.630 ;
        RECT 131.680 205.150 134.420 205.220 ;
        RECT 131.550 205.050 134.420 205.150 ;
        RECT 131.550 203.640 131.850 205.050 ;
        RECT 132.190 204.180 132.360 204.510 ;
        RECT 132.530 204.480 133.570 204.650 ;
        RECT 132.530 204.040 133.570 204.210 ;
        RECT 133.740 204.180 133.910 204.510 ;
        RECT 134.250 203.640 134.420 205.050 ;
        RECT 131.550 203.500 134.420 203.640 ;
        RECT 131.680 203.470 134.420 203.500 ;
        RECT 134.980 205.180 137.810 205.230 ;
        RECT 153.730 205.220 156.470 205.290 ;
        RECT 134.980 205.060 137.930 205.180 ;
        RECT 134.980 203.650 135.150 205.060 ;
        RECT 135.490 204.190 135.660 204.520 ;
        RECT 135.875 204.490 136.915 204.660 ;
        RECT 135.875 204.050 136.915 204.220 ;
        RECT 137.130 204.190 137.300 204.520 ;
        RECT 137.640 203.650 137.930 205.060 ;
        RECT 134.980 203.530 137.930 203.650 ;
        RECT 153.600 205.120 156.470 205.220 ;
        RECT 153.600 203.710 153.900 205.120 ;
        RECT 154.240 204.250 154.410 204.580 ;
        RECT 154.580 204.550 155.620 204.720 ;
        RECT 154.580 204.110 155.620 204.280 ;
        RECT 155.790 204.250 155.960 204.580 ;
        RECT 156.300 203.710 156.470 205.120 ;
        RECT 153.600 203.570 156.470 203.710 ;
        RECT 153.730 203.540 156.470 203.570 ;
        RECT 157.030 205.250 159.860 205.300 ;
        RECT 157.030 205.130 159.980 205.250 ;
        RECT 157.030 203.720 157.200 205.130 ;
        RECT 157.540 204.260 157.710 204.590 ;
        RECT 157.925 204.560 158.965 204.730 ;
        RECT 157.925 204.120 158.965 204.290 ;
        RECT 159.180 204.260 159.350 204.590 ;
        RECT 159.690 203.720 159.980 205.130 ;
        RECT 157.030 203.600 159.980 203.720 ;
        RECT 157.030 203.550 159.860 203.600 ;
        RECT 134.980 203.480 137.810 203.530 ;
        RECT 131.680 203.060 134.420 203.130 ;
        RECT 131.550 202.960 134.420 203.060 ;
        RECT 131.550 201.550 131.850 202.960 ;
        RECT 132.190 202.090 132.360 202.420 ;
        RECT 132.530 202.390 133.570 202.560 ;
        RECT 132.530 201.950 133.570 202.120 ;
        RECT 133.740 202.090 133.910 202.420 ;
        RECT 134.250 201.550 134.420 202.960 ;
        RECT 131.550 201.410 134.420 201.550 ;
        RECT 131.680 201.380 134.420 201.410 ;
        RECT 134.980 203.090 137.810 203.140 ;
        RECT 153.730 203.120 156.470 203.190 ;
        RECT 134.980 202.970 137.930 203.090 ;
        RECT 134.980 201.560 135.150 202.970 ;
        RECT 135.490 202.100 135.660 202.430 ;
        RECT 135.875 202.400 136.915 202.570 ;
        RECT 135.875 201.960 136.915 202.130 ;
        RECT 137.130 202.100 137.300 202.430 ;
        RECT 137.640 201.560 137.930 202.970 ;
        RECT 134.980 201.440 137.930 201.560 ;
        RECT 153.600 203.020 156.470 203.120 ;
        RECT 153.600 201.610 153.900 203.020 ;
        RECT 154.240 202.150 154.410 202.480 ;
        RECT 154.580 202.450 155.620 202.620 ;
        RECT 154.580 202.010 155.620 202.180 ;
        RECT 155.790 202.150 155.960 202.480 ;
        RECT 156.300 201.610 156.470 203.020 ;
        RECT 153.600 201.470 156.470 201.610 ;
        RECT 153.730 201.440 156.470 201.470 ;
        RECT 157.030 203.150 159.860 203.200 ;
        RECT 157.030 203.030 159.980 203.150 ;
        RECT 157.030 201.620 157.200 203.030 ;
        RECT 157.540 202.160 157.710 202.490 ;
        RECT 157.925 202.460 158.965 202.630 ;
        RECT 157.925 202.020 158.965 202.190 ;
        RECT 159.180 202.160 159.350 202.490 ;
        RECT 159.690 201.620 159.980 203.030 ;
        RECT 157.030 201.500 159.980 201.620 ;
        RECT 157.030 201.450 159.860 201.500 ;
        RECT 134.980 201.390 137.810 201.440 ;
        RECT 131.680 200.960 134.420 201.030 ;
        RECT 131.550 200.860 134.420 200.960 ;
        RECT 131.550 199.450 131.850 200.860 ;
        RECT 132.190 199.990 132.360 200.320 ;
        RECT 132.530 200.290 133.570 200.460 ;
        RECT 132.530 199.850 133.570 200.020 ;
        RECT 133.740 199.990 133.910 200.320 ;
        RECT 134.250 199.450 134.420 200.860 ;
        RECT 131.550 199.310 134.420 199.450 ;
        RECT 131.680 199.280 134.420 199.310 ;
        RECT 134.980 200.990 137.810 201.040 ;
        RECT 153.730 201.020 156.470 201.090 ;
        RECT 134.980 200.870 137.930 200.990 ;
        RECT 134.980 199.460 135.150 200.870 ;
        RECT 135.490 200.000 135.660 200.330 ;
        RECT 135.875 200.300 136.915 200.470 ;
        RECT 135.875 199.860 136.915 200.030 ;
        RECT 137.130 200.000 137.300 200.330 ;
        RECT 137.640 199.460 137.930 200.870 ;
        RECT 134.980 199.340 137.930 199.460 ;
        RECT 153.600 200.920 156.470 201.020 ;
        RECT 153.600 199.510 153.900 200.920 ;
        RECT 154.240 200.050 154.410 200.380 ;
        RECT 154.580 200.350 155.620 200.520 ;
        RECT 154.580 199.910 155.620 200.080 ;
        RECT 155.790 200.050 155.960 200.380 ;
        RECT 156.300 199.510 156.470 200.920 ;
        RECT 153.600 199.370 156.470 199.510 ;
        RECT 153.730 199.340 156.470 199.370 ;
        RECT 157.030 201.050 159.860 201.100 ;
        RECT 157.030 200.930 159.980 201.050 ;
        RECT 157.030 199.520 157.200 200.930 ;
        RECT 157.540 200.060 157.710 200.390 ;
        RECT 157.925 200.360 158.965 200.530 ;
        RECT 157.925 199.920 158.965 200.090 ;
        RECT 159.180 200.060 159.350 200.390 ;
        RECT 159.690 199.520 159.980 200.930 ;
        RECT 157.030 199.400 159.980 199.520 ;
        RECT 157.030 199.350 159.860 199.400 ;
        RECT 134.980 199.290 137.810 199.340 ;
        RECT 131.680 198.870 134.420 198.940 ;
        RECT 131.550 198.770 134.420 198.870 ;
        RECT 131.550 197.360 131.850 198.770 ;
        RECT 132.190 197.900 132.360 198.230 ;
        RECT 132.530 198.200 133.570 198.370 ;
        RECT 132.530 197.760 133.570 197.930 ;
        RECT 133.740 197.900 133.910 198.230 ;
        RECT 134.250 197.360 134.420 198.770 ;
        RECT 131.550 197.220 134.420 197.360 ;
        RECT 131.680 197.190 134.420 197.220 ;
        RECT 134.980 198.900 137.810 198.950 ;
        RECT 153.730 198.920 156.470 198.990 ;
        RECT 134.980 198.780 137.930 198.900 ;
        RECT 134.980 197.370 135.150 198.780 ;
        RECT 135.490 197.910 135.660 198.240 ;
        RECT 135.875 198.210 136.915 198.380 ;
        RECT 135.875 197.770 136.915 197.940 ;
        RECT 137.130 197.910 137.300 198.240 ;
        RECT 137.640 197.370 137.930 198.780 ;
        RECT 134.980 197.250 137.930 197.370 ;
        RECT 153.600 198.820 156.470 198.920 ;
        RECT 153.600 197.410 153.900 198.820 ;
        RECT 154.240 197.950 154.410 198.280 ;
        RECT 154.580 198.250 155.620 198.420 ;
        RECT 154.580 197.810 155.620 197.980 ;
        RECT 155.790 197.950 155.960 198.280 ;
        RECT 156.300 197.410 156.470 198.820 ;
        RECT 153.600 197.270 156.470 197.410 ;
        RECT 134.980 197.200 137.810 197.250 ;
        RECT 153.730 197.240 156.470 197.270 ;
        RECT 157.030 198.950 159.860 199.000 ;
        RECT 157.030 198.830 159.980 198.950 ;
        RECT 157.030 197.420 157.200 198.830 ;
        RECT 157.540 197.960 157.710 198.290 ;
        RECT 157.925 198.260 158.965 198.430 ;
        RECT 157.925 197.820 158.965 197.990 ;
        RECT 159.180 197.960 159.350 198.290 ;
        RECT 159.690 197.420 159.980 198.830 ;
        RECT 157.030 197.300 159.980 197.420 ;
        RECT 157.030 197.250 159.860 197.300 ;
        RECT 131.680 196.770 134.420 196.840 ;
        RECT 131.550 196.670 134.420 196.770 ;
        RECT 131.550 195.260 131.850 196.670 ;
        RECT 132.190 195.800 132.360 196.130 ;
        RECT 132.530 196.100 133.570 196.270 ;
        RECT 132.530 195.660 133.570 195.830 ;
        RECT 133.740 195.800 133.910 196.130 ;
        RECT 134.250 195.260 134.420 196.670 ;
        RECT 131.550 195.120 134.420 195.260 ;
        RECT 131.680 195.090 134.420 195.120 ;
        RECT 134.980 196.800 137.810 196.850 ;
        RECT 153.730 196.820 156.470 196.890 ;
        RECT 134.980 196.680 137.930 196.800 ;
        RECT 134.980 195.270 135.150 196.680 ;
        RECT 135.490 195.810 135.660 196.140 ;
        RECT 135.875 196.110 136.915 196.280 ;
        RECT 135.875 195.670 136.915 195.840 ;
        RECT 137.130 195.810 137.300 196.140 ;
        RECT 137.640 195.270 137.930 196.680 ;
        RECT 134.980 195.150 137.930 195.270 ;
        RECT 153.600 196.720 156.470 196.820 ;
        RECT 153.600 195.310 153.900 196.720 ;
        RECT 154.240 195.850 154.410 196.180 ;
        RECT 154.580 196.150 155.620 196.320 ;
        RECT 154.580 195.710 155.620 195.880 ;
        RECT 155.790 195.850 155.960 196.180 ;
        RECT 156.300 195.310 156.470 196.720 ;
        RECT 153.600 195.170 156.470 195.310 ;
        RECT 134.980 195.100 137.810 195.150 ;
        RECT 153.730 195.140 156.470 195.170 ;
        RECT 157.030 196.850 159.860 196.900 ;
        RECT 157.030 196.730 159.980 196.850 ;
        RECT 157.030 195.320 157.200 196.730 ;
        RECT 157.540 195.860 157.710 196.190 ;
        RECT 157.925 196.160 158.965 196.330 ;
        RECT 157.925 195.720 158.965 195.890 ;
        RECT 159.180 195.860 159.350 196.190 ;
        RECT 159.690 195.320 159.980 196.730 ;
        RECT 157.030 195.200 159.980 195.320 ;
        RECT 157.030 195.150 159.860 195.200 ;
        RECT 131.680 194.670 134.420 194.740 ;
        RECT 131.550 194.570 134.420 194.670 ;
        RECT 131.550 193.160 131.850 194.570 ;
        RECT 132.190 193.700 132.360 194.030 ;
        RECT 132.530 194.000 133.570 194.170 ;
        RECT 132.530 193.560 133.570 193.730 ;
        RECT 133.740 193.700 133.910 194.030 ;
        RECT 134.250 193.160 134.420 194.570 ;
        RECT 131.550 193.020 134.420 193.160 ;
        RECT 131.680 192.990 134.420 193.020 ;
        RECT 134.980 194.700 137.810 194.750 ;
        RECT 153.730 194.720 156.470 194.790 ;
        RECT 134.980 194.580 137.930 194.700 ;
        RECT 134.980 193.170 135.150 194.580 ;
        RECT 135.490 193.710 135.660 194.040 ;
        RECT 135.875 194.010 136.915 194.180 ;
        RECT 135.875 193.570 136.915 193.740 ;
        RECT 137.130 193.710 137.300 194.040 ;
        RECT 137.640 193.170 137.930 194.580 ;
        RECT 134.980 193.050 137.930 193.170 ;
        RECT 153.600 194.620 156.470 194.720 ;
        RECT 153.600 193.210 153.900 194.620 ;
        RECT 154.240 193.750 154.410 194.080 ;
        RECT 154.580 194.050 155.620 194.220 ;
        RECT 154.580 193.610 155.620 193.780 ;
        RECT 155.790 193.750 155.960 194.080 ;
        RECT 156.300 193.210 156.470 194.620 ;
        RECT 153.600 193.070 156.470 193.210 ;
        RECT 134.980 193.000 137.810 193.050 ;
        RECT 153.730 193.040 156.470 193.070 ;
        RECT 157.030 194.750 159.860 194.800 ;
        RECT 157.030 194.630 159.980 194.750 ;
        RECT 157.030 193.220 157.200 194.630 ;
        RECT 157.540 193.760 157.710 194.090 ;
        RECT 157.925 194.060 158.965 194.230 ;
        RECT 157.925 193.620 158.965 193.790 ;
        RECT 159.180 193.760 159.350 194.090 ;
        RECT 159.690 193.220 159.980 194.630 ;
        RECT 157.030 193.100 159.980 193.220 ;
        RECT 157.030 193.050 159.860 193.100 ;
        RECT 131.680 192.570 134.420 192.640 ;
        RECT 131.550 192.470 134.420 192.570 ;
        RECT 131.550 191.060 131.850 192.470 ;
        RECT 132.190 191.600 132.360 191.930 ;
        RECT 132.530 191.900 133.570 192.070 ;
        RECT 132.530 191.460 133.570 191.630 ;
        RECT 133.740 191.600 133.910 191.930 ;
        RECT 134.250 191.060 134.420 192.470 ;
        RECT 131.550 190.920 134.420 191.060 ;
        RECT 131.680 190.890 134.420 190.920 ;
        RECT 134.980 192.600 137.810 192.650 ;
        RECT 153.730 192.620 156.470 192.690 ;
        RECT 134.980 192.480 137.930 192.600 ;
        RECT 134.980 191.070 135.150 192.480 ;
        RECT 135.490 191.610 135.660 191.940 ;
        RECT 135.875 191.910 136.915 192.080 ;
        RECT 135.875 191.470 136.915 191.640 ;
        RECT 137.130 191.610 137.300 191.940 ;
        RECT 137.640 191.070 137.930 192.480 ;
        RECT 134.980 190.950 137.930 191.070 ;
        RECT 153.600 192.520 156.470 192.620 ;
        RECT 153.600 191.110 153.900 192.520 ;
        RECT 154.240 191.650 154.410 191.980 ;
        RECT 154.580 191.950 155.620 192.120 ;
        RECT 154.580 191.510 155.620 191.680 ;
        RECT 155.790 191.650 155.960 191.980 ;
        RECT 156.300 191.110 156.470 192.520 ;
        RECT 153.600 190.970 156.470 191.110 ;
        RECT 134.980 190.900 137.810 190.950 ;
        RECT 153.730 190.940 156.470 190.970 ;
        RECT 157.030 192.650 159.860 192.700 ;
        RECT 157.030 192.530 159.980 192.650 ;
        RECT 157.030 191.120 157.200 192.530 ;
        RECT 157.540 191.660 157.710 191.990 ;
        RECT 157.925 191.960 158.965 192.130 ;
        RECT 157.925 191.520 158.965 191.690 ;
        RECT 159.180 191.660 159.350 191.990 ;
        RECT 159.690 191.120 159.980 192.530 ;
        RECT 157.030 191.000 159.980 191.120 ;
        RECT 157.030 190.950 159.860 191.000 ;
        RECT 131.680 190.470 134.420 190.540 ;
        RECT 131.550 190.370 134.420 190.470 ;
        RECT 131.550 188.960 131.850 190.370 ;
        RECT 132.190 189.500 132.360 189.830 ;
        RECT 132.530 189.800 133.570 189.970 ;
        RECT 132.530 189.360 133.570 189.530 ;
        RECT 133.740 189.500 133.910 189.830 ;
        RECT 134.250 188.960 134.420 190.370 ;
        RECT 131.550 188.820 134.420 188.960 ;
        RECT 131.680 188.790 134.420 188.820 ;
        RECT 134.980 190.500 137.810 190.550 ;
        RECT 153.730 190.520 156.470 190.590 ;
        RECT 134.980 190.380 137.930 190.500 ;
        RECT 134.980 188.970 135.150 190.380 ;
        RECT 135.490 189.510 135.660 189.840 ;
        RECT 135.875 189.810 136.915 189.980 ;
        RECT 135.875 189.370 136.915 189.540 ;
        RECT 137.130 189.510 137.300 189.840 ;
        RECT 137.640 188.970 137.930 190.380 ;
        RECT 134.980 188.850 137.930 188.970 ;
        RECT 153.600 190.420 156.470 190.520 ;
        RECT 153.600 189.010 153.900 190.420 ;
        RECT 154.240 189.550 154.410 189.880 ;
        RECT 154.580 189.850 155.620 190.020 ;
        RECT 154.580 189.410 155.620 189.580 ;
        RECT 155.790 189.550 155.960 189.880 ;
        RECT 156.300 189.010 156.470 190.420 ;
        RECT 153.600 188.870 156.470 189.010 ;
        RECT 134.980 188.800 137.810 188.850 ;
        RECT 153.730 188.840 156.470 188.870 ;
        RECT 157.030 190.550 159.860 190.600 ;
        RECT 157.030 190.430 159.980 190.550 ;
        RECT 157.030 189.020 157.200 190.430 ;
        RECT 157.540 189.560 157.710 189.890 ;
        RECT 157.925 189.860 158.965 190.030 ;
        RECT 157.925 189.420 158.965 189.590 ;
        RECT 159.180 189.560 159.350 189.890 ;
        RECT 159.690 189.020 159.980 190.430 ;
        RECT 157.030 188.900 159.980 189.020 ;
        RECT 157.030 188.850 159.860 188.900 ;
        RECT 131.680 188.370 134.420 188.440 ;
        RECT 131.550 188.270 134.420 188.370 ;
        RECT 131.550 186.860 131.850 188.270 ;
        RECT 132.190 187.400 132.360 187.730 ;
        RECT 132.530 187.700 133.570 187.870 ;
        RECT 132.530 187.260 133.570 187.430 ;
        RECT 133.740 187.400 133.910 187.730 ;
        RECT 134.250 186.860 134.420 188.270 ;
        RECT 131.550 186.720 134.420 186.860 ;
        RECT 131.680 186.690 134.420 186.720 ;
        RECT 134.980 188.400 137.810 188.450 ;
        RECT 153.730 188.420 156.470 188.490 ;
        RECT 134.980 188.280 137.930 188.400 ;
        RECT 134.980 186.870 135.150 188.280 ;
        RECT 135.490 187.410 135.660 187.740 ;
        RECT 135.875 187.710 136.915 187.880 ;
        RECT 135.875 187.270 136.915 187.440 ;
        RECT 137.130 187.410 137.300 187.740 ;
        RECT 137.640 186.870 137.930 188.280 ;
        RECT 134.980 186.750 137.930 186.870 ;
        RECT 153.600 188.320 156.470 188.420 ;
        RECT 153.600 186.910 153.900 188.320 ;
        RECT 154.240 187.450 154.410 187.780 ;
        RECT 154.580 187.750 155.620 187.920 ;
        RECT 154.580 187.310 155.620 187.480 ;
        RECT 155.790 187.450 155.960 187.780 ;
        RECT 156.300 186.910 156.470 188.320 ;
        RECT 153.600 186.770 156.470 186.910 ;
        RECT 134.980 186.700 137.810 186.750 ;
        RECT 153.730 186.740 156.470 186.770 ;
        RECT 157.030 188.450 159.860 188.500 ;
        RECT 157.030 188.330 159.980 188.450 ;
        RECT 157.030 186.920 157.200 188.330 ;
        RECT 157.540 187.460 157.710 187.790 ;
        RECT 157.925 187.760 158.965 187.930 ;
        RECT 157.925 187.320 158.965 187.490 ;
        RECT 159.180 187.460 159.350 187.790 ;
        RECT 159.690 186.920 159.980 188.330 ;
        RECT 157.030 186.800 159.980 186.920 ;
        RECT 157.030 186.750 159.860 186.800 ;
        RECT 131.680 186.270 134.420 186.340 ;
        RECT 131.550 186.170 134.420 186.270 ;
        RECT 131.550 184.760 131.850 186.170 ;
        RECT 132.190 185.300 132.360 185.630 ;
        RECT 132.530 185.600 133.570 185.770 ;
        RECT 132.530 185.160 133.570 185.330 ;
        RECT 133.740 185.300 133.910 185.630 ;
        RECT 134.250 184.760 134.420 186.170 ;
        RECT 131.550 184.620 134.420 184.760 ;
        RECT 131.680 184.590 134.420 184.620 ;
        RECT 134.980 186.300 137.810 186.350 ;
        RECT 153.730 186.320 156.470 186.390 ;
        RECT 134.980 186.180 137.930 186.300 ;
        RECT 134.980 184.770 135.150 186.180 ;
        RECT 135.490 185.310 135.660 185.640 ;
        RECT 135.875 185.610 136.915 185.780 ;
        RECT 135.875 185.170 136.915 185.340 ;
        RECT 137.130 185.310 137.300 185.640 ;
        RECT 137.640 184.770 137.930 186.180 ;
        RECT 134.980 184.650 137.930 184.770 ;
        RECT 153.600 186.220 156.470 186.320 ;
        RECT 153.600 184.810 153.900 186.220 ;
        RECT 154.240 185.350 154.410 185.680 ;
        RECT 154.580 185.650 155.620 185.820 ;
        RECT 154.580 185.210 155.620 185.380 ;
        RECT 155.790 185.350 155.960 185.680 ;
        RECT 156.300 184.810 156.470 186.220 ;
        RECT 153.600 184.670 156.470 184.810 ;
        RECT 134.980 184.600 137.810 184.650 ;
        RECT 153.730 184.640 156.470 184.670 ;
        RECT 157.030 186.350 159.860 186.400 ;
        RECT 157.030 186.230 159.980 186.350 ;
        RECT 157.030 184.820 157.200 186.230 ;
        RECT 157.540 185.360 157.710 185.690 ;
        RECT 157.925 185.660 158.965 185.830 ;
        RECT 157.925 185.220 158.965 185.390 ;
        RECT 159.180 185.360 159.350 185.690 ;
        RECT 159.690 184.820 159.980 186.230 ;
        RECT 157.030 184.700 159.980 184.820 ;
        RECT 157.030 184.650 159.860 184.700 ;
        RECT 131.680 184.170 134.420 184.240 ;
        RECT 131.550 184.070 134.420 184.170 ;
        RECT 131.550 182.660 131.850 184.070 ;
        RECT 132.190 183.200 132.360 183.530 ;
        RECT 132.530 183.500 133.570 183.670 ;
        RECT 132.530 183.060 133.570 183.230 ;
        RECT 133.740 183.200 133.910 183.530 ;
        RECT 134.250 182.660 134.420 184.070 ;
        RECT 131.550 182.520 134.420 182.660 ;
        RECT 131.680 182.490 134.420 182.520 ;
        RECT 134.980 184.200 137.810 184.250 ;
        RECT 153.730 184.220 156.470 184.290 ;
        RECT 134.980 184.080 137.930 184.200 ;
        RECT 134.980 182.670 135.150 184.080 ;
        RECT 135.490 183.210 135.660 183.540 ;
        RECT 135.875 183.510 136.915 183.680 ;
        RECT 135.875 183.070 136.915 183.240 ;
        RECT 137.130 183.210 137.300 183.540 ;
        RECT 137.640 182.670 137.930 184.080 ;
        RECT 134.980 182.550 137.930 182.670 ;
        RECT 153.600 184.120 156.470 184.220 ;
        RECT 153.600 182.710 153.900 184.120 ;
        RECT 154.240 183.250 154.410 183.580 ;
        RECT 154.580 183.550 155.620 183.720 ;
        RECT 154.580 183.110 155.620 183.280 ;
        RECT 155.790 183.250 155.960 183.580 ;
        RECT 156.300 182.710 156.470 184.120 ;
        RECT 153.600 182.570 156.470 182.710 ;
        RECT 134.980 182.500 137.810 182.550 ;
        RECT 153.730 182.540 156.470 182.570 ;
        RECT 157.030 184.250 159.860 184.300 ;
        RECT 157.030 184.130 159.980 184.250 ;
        RECT 157.030 182.720 157.200 184.130 ;
        RECT 157.540 183.260 157.710 183.590 ;
        RECT 157.925 183.560 158.965 183.730 ;
        RECT 157.925 183.120 158.965 183.290 ;
        RECT 159.180 183.260 159.350 183.590 ;
        RECT 159.690 182.720 159.980 184.130 ;
        RECT 157.030 182.600 159.980 182.720 ;
        RECT 157.030 182.550 159.860 182.600 ;
        RECT 131.680 182.070 134.420 182.140 ;
        RECT 131.550 181.970 134.420 182.070 ;
        RECT 131.550 180.560 131.850 181.970 ;
        RECT 132.190 181.100 132.360 181.430 ;
        RECT 132.530 181.400 133.570 181.570 ;
        RECT 132.530 180.960 133.570 181.130 ;
        RECT 133.740 181.100 133.910 181.430 ;
        RECT 134.250 180.560 134.420 181.970 ;
        RECT 131.550 180.420 134.420 180.560 ;
        RECT 131.680 180.390 134.420 180.420 ;
        RECT 134.980 182.100 137.810 182.150 ;
        RECT 153.730 182.120 156.470 182.190 ;
        RECT 134.980 181.980 137.930 182.100 ;
        RECT 134.980 180.570 135.150 181.980 ;
        RECT 135.490 181.110 135.660 181.440 ;
        RECT 135.875 181.410 136.915 181.580 ;
        RECT 135.875 180.970 136.915 181.140 ;
        RECT 137.130 181.110 137.300 181.440 ;
        RECT 137.640 180.570 137.930 181.980 ;
        RECT 134.980 180.450 137.930 180.570 ;
        RECT 153.600 182.020 156.470 182.120 ;
        RECT 153.600 180.610 153.900 182.020 ;
        RECT 154.240 181.150 154.410 181.480 ;
        RECT 154.580 181.450 155.620 181.620 ;
        RECT 154.580 181.010 155.620 181.180 ;
        RECT 155.790 181.150 155.960 181.480 ;
        RECT 156.300 180.610 156.470 182.020 ;
        RECT 153.600 180.470 156.470 180.610 ;
        RECT 134.980 180.400 137.810 180.450 ;
        RECT 153.730 180.440 156.470 180.470 ;
        RECT 157.030 182.150 159.860 182.200 ;
        RECT 157.030 182.030 159.980 182.150 ;
        RECT 157.030 180.620 157.200 182.030 ;
        RECT 157.540 181.160 157.710 181.490 ;
        RECT 157.925 181.460 158.965 181.630 ;
        RECT 157.925 181.020 158.965 181.190 ;
        RECT 159.180 181.160 159.350 181.490 ;
        RECT 159.690 180.620 159.980 182.030 ;
        RECT 157.030 180.500 159.980 180.620 ;
        RECT 157.030 180.450 159.860 180.500 ;
        RECT 131.680 179.980 134.420 180.050 ;
        RECT 131.550 179.880 134.420 179.980 ;
        RECT 131.550 178.470 131.850 179.880 ;
        RECT 132.190 179.010 132.360 179.340 ;
        RECT 132.530 179.310 133.570 179.480 ;
        RECT 132.530 178.870 133.570 179.040 ;
        RECT 133.740 179.010 133.910 179.340 ;
        RECT 134.250 178.470 134.420 179.880 ;
        RECT 131.550 178.330 134.420 178.470 ;
        RECT 131.680 178.300 134.420 178.330 ;
        RECT 134.980 180.010 137.810 180.060 ;
        RECT 153.730 180.020 156.470 180.090 ;
        RECT 134.980 179.890 137.930 180.010 ;
        RECT 134.980 178.480 135.150 179.890 ;
        RECT 135.490 179.020 135.660 179.350 ;
        RECT 135.875 179.320 136.915 179.490 ;
        RECT 135.875 178.880 136.915 179.050 ;
        RECT 137.130 179.020 137.300 179.350 ;
        RECT 137.640 178.480 137.930 179.890 ;
        RECT 134.980 178.360 137.930 178.480 ;
        RECT 153.600 179.920 156.470 180.020 ;
        RECT 153.600 178.510 153.900 179.920 ;
        RECT 154.240 179.050 154.410 179.380 ;
        RECT 154.580 179.350 155.620 179.520 ;
        RECT 154.580 178.910 155.620 179.080 ;
        RECT 155.790 179.050 155.960 179.380 ;
        RECT 156.300 178.510 156.470 179.920 ;
        RECT 153.600 178.370 156.470 178.510 ;
        RECT 134.980 178.310 137.810 178.360 ;
        RECT 153.730 178.340 156.470 178.370 ;
        RECT 157.030 180.050 159.860 180.100 ;
        RECT 157.030 179.930 159.980 180.050 ;
        RECT 157.030 178.520 157.200 179.930 ;
        RECT 157.540 179.060 157.710 179.390 ;
        RECT 157.925 179.360 158.965 179.530 ;
        RECT 157.925 178.920 158.965 179.090 ;
        RECT 159.180 179.060 159.350 179.390 ;
        RECT 159.690 178.520 159.980 179.930 ;
        RECT 157.030 178.400 159.980 178.520 ;
        RECT 157.030 178.350 159.860 178.400 ;
        RECT 131.680 177.890 134.420 177.960 ;
        RECT 131.550 177.790 134.420 177.890 ;
        RECT 131.550 176.380 131.850 177.790 ;
        RECT 132.190 176.920 132.360 177.250 ;
        RECT 132.530 177.220 133.570 177.390 ;
        RECT 132.530 176.780 133.570 176.950 ;
        RECT 133.740 176.920 133.910 177.250 ;
        RECT 134.250 176.380 134.420 177.790 ;
        RECT 131.550 176.240 134.420 176.380 ;
        RECT 131.680 176.210 134.420 176.240 ;
        RECT 134.980 177.920 137.810 177.970 ;
        RECT 153.730 177.920 156.470 177.990 ;
        RECT 134.980 177.800 137.930 177.920 ;
        RECT 134.980 176.390 135.150 177.800 ;
        RECT 135.490 176.930 135.660 177.260 ;
        RECT 135.875 177.230 136.915 177.400 ;
        RECT 135.875 176.790 136.915 176.960 ;
        RECT 137.130 176.930 137.300 177.260 ;
        RECT 137.640 176.390 137.930 177.800 ;
        RECT 134.980 176.270 137.930 176.390 ;
        RECT 153.600 177.820 156.470 177.920 ;
        RECT 153.600 176.410 153.900 177.820 ;
        RECT 154.240 176.950 154.410 177.280 ;
        RECT 154.580 177.250 155.620 177.420 ;
        RECT 154.580 176.810 155.620 176.980 ;
        RECT 155.790 176.950 155.960 177.280 ;
        RECT 156.300 176.410 156.470 177.820 ;
        RECT 153.600 176.270 156.470 176.410 ;
        RECT 134.980 176.220 137.810 176.270 ;
        RECT 153.730 176.240 156.470 176.270 ;
        RECT 157.030 177.950 159.860 178.000 ;
        RECT 157.030 177.830 159.980 177.950 ;
        RECT 157.030 176.420 157.200 177.830 ;
        RECT 157.540 176.960 157.710 177.290 ;
        RECT 157.925 177.260 158.965 177.430 ;
        RECT 157.925 176.820 158.965 176.990 ;
        RECT 159.180 176.960 159.350 177.290 ;
        RECT 159.690 176.420 159.980 177.830 ;
        RECT 157.030 176.300 159.980 176.420 ;
        RECT 157.030 176.250 159.860 176.300 ;
        RECT 131.680 175.790 134.420 175.860 ;
        RECT 131.550 175.690 134.420 175.790 ;
        RECT 131.550 174.280 131.850 175.690 ;
        RECT 132.190 174.820 132.360 175.150 ;
        RECT 132.530 175.120 133.570 175.290 ;
        RECT 132.530 174.680 133.570 174.850 ;
        RECT 133.740 174.820 133.910 175.150 ;
        RECT 134.250 174.280 134.420 175.690 ;
        RECT 131.550 174.140 134.420 174.280 ;
        RECT 131.680 174.110 134.420 174.140 ;
        RECT 134.980 175.820 137.810 175.870 ;
        RECT 153.730 175.820 156.470 175.890 ;
        RECT 134.980 175.700 137.930 175.820 ;
        RECT 134.980 174.290 135.150 175.700 ;
        RECT 135.490 174.830 135.660 175.160 ;
        RECT 135.875 175.130 136.915 175.300 ;
        RECT 135.875 174.690 136.915 174.860 ;
        RECT 137.130 174.830 137.300 175.160 ;
        RECT 137.640 174.290 137.930 175.700 ;
        RECT 134.980 174.170 137.930 174.290 ;
        RECT 153.600 175.720 156.470 175.820 ;
        RECT 153.600 174.310 153.900 175.720 ;
        RECT 154.240 174.850 154.410 175.180 ;
        RECT 154.580 175.150 155.620 175.320 ;
        RECT 154.580 174.710 155.620 174.880 ;
        RECT 155.790 174.850 155.960 175.180 ;
        RECT 156.300 174.310 156.470 175.720 ;
        RECT 153.600 174.170 156.470 174.310 ;
        RECT 134.980 174.120 137.810 174.170 ;
        RECT 153.730 174.140 156.470 174.170 ;
        RECT 157.030 175.850 159.860 175.900 ;
        RECT 157.030 175.730 159.980 175.850 ;
        RECT 157.030 174.320 157.200 175.730 ;
        RECT 157.540 174.860 157.710 175.190 ;
        RECT 157.925 175.160 158.965 175.330 ;
        RECT 157.925 174.720 158.965 174.890 ;
        RECT 159.180 174.860 159.350 175.190 ;
        RECT 159.690 174.320 159.980 175.730 ;
        RECT 157.030 174.200 159.980 174.320 ;
        RECT 157.030 174.150 159.860 174.200 ;
        RECT 131.680 173.700 134.420 173.770 ;
        RECT 131.550 173.600 134.420 173.700 ;
        RECT 131.550 172.190 131.850 173.600 ;
        RECT 132.190 172.730 132.360 173.060 ;
        RECT 132.530 173.030 133.570 173.200 ;
        RECT 132.530 172.590 133.570 172.760 ;
        RECT 133.740 172.730 133.910 173.060 ;
        RECT 134.250 172.190 134.420 173.600 ;
        RECT 131.550 172.050 134.420 172.190 ;
        RECT 131.680 172.020 134.420 172.050 ;
        RECT 134.980 173.730 137.810 173.780 ;
        RECT 134.980 173.610 137.930 173.730 ;
        RECT 153.730 173.720 156.470 173.790 ;
        RECT 134.980 172.200 135.150 173.610 ;
        RECT 135.490 172.740 135.660 173.070 ;
        RECT 135.875 173.040 136.915 173.210 ;
        RECT 135.875 172.600 136.915 172.770 ;
        RECT 137.130 172.740 137.300 173.070 ;
        RECT 137.640 172.200 137.930 173.610 ;
        RECT 134.980 172.080 137.930 172.200 ;
        RECT 153.600 173.620 156.470 173.720 ;
        RECT 153.600 172.210 153.900 173.620 ;
        RECT 154.240 172.750 154.410 173.080 ;
        RECT 154.580 173.050 155.620 173.220 ;
        RECT 154.580 172.610 155.620 172.780 ;
        RECT 155.790 172.750 155.960 173.080 ;
        RECT 156.300 172.210 156.470 173.620 ;
        RECT 134.980 172.030 137.810 172.080 ;
        RECT 153.600 172.070 156.470 172.210 ;
        RECT 153.730 172.040 156.470 172.070 ;
        RECT 157.030 173.750 159.860 173.800 ;
        RECT 157.030 173.630 159.980 173.750 ;
        RECT 157.030 172.220 157.200 173.630 ;
        RECT 157.540 172.760 157.710 173.090 ;
        RECT 157.925 173.060 158.965 173.230 ;
        RECT 157.925 172.620 158.965 172.790 ;
        RECT 159.180 172.760 159.350 173.090 ;
        RECT 159.690 172.220 159.980 173.630 ;
        RECT 157.030 172.100 159.980 172.220 ;
        RECT 157.030 172.050 159.860 172.100 ;
        RECT 131.680 171.610 134.420 171.680 ;
        RECT 131.550 171.510 134.420 171.610 ;
        RECT 131.550 170.100 131.850 171.510 ;
        RECT 132.190 170.640 132.360 170.970 ;
        RECT 132.530 170.940 133.570 171.110 ;
        RECT 132.530 170.500 133.570 170.670 ;
        RECT 133.740 170.640 133.910 170.970 ;
        RECT 134.250 170.100 134.420 171.510 ;
        RECT 131.550 169.960 134.420 170.100 ;
        RECT 131.680 169.930 134.420 169.960 ;
        RECT 134.980 171.640 137.810 171.690 ;
        RECT 134.980 171.520 137.930 171.640 ;
        RECT 153.730 171.620 156.470 171.690 ;
        RECT 134.980 170.110 135.150 171.520 ;
        RECT 135.490 170.650 135.660 170.980 ;
        RECT 135.875 170.950 136.915 171.120 ;
        RECT 135.875 170.510 136.915 170.680 ;
        RECT 137.130 170.650 137.300 170.980 ;
        RECT 137.640 170.110 137.930 171.520 ;
        RECT 134.980 169.990 137.930 170.110 ;
        RECT 153.600 171.520 156.470 171.620 ;
        RECT 153.600 170.110 153.900 171.520 ;
        RECT 154.240 170.650 154.410 170.980 ;
        RECT 154.580 170.950 155.620 171.120 ;
        RECT 154.580 170.510 155.620 170.680 ;
        RECT 155.790 170.650 155.960 170.980 ;
        RECT 156.300 170.110 156.470 171.520 ;
        RECT 134.980 169.940 137.810 169.990 ;
        RECT 153.600 169.970 156.470 170.110 ;
        RECT 153.730 169.940 156.470 169.970 ;
        RECT 157.030 171.650 159.860 171.700 ;
        RECT 157.030 171.530 159.980 171.650 ;
        RECT 157.030 170.120 157.200 171.530 ;
        RECT 157.540 170.660 157.710 170.990 ;
        RECT 157.925 170.960 158.965 171.130 ;
        RECT 157.925 170.520 158.965 170.690 ;
        RECT 159.180 170.660 159.350 170.990 ;
        RECT 159.690 170.120 159.980 171.530 ;
        RECT 157.030 170.000 159.980 170.120 ;
        RECT 157.030 169.950 159.860 170.000 ;
        RECT 131.680 169.510 134.420 169.580 ;
        RECT 131.550 169.410 134.420 169.510 ;
        RECT 131.550 168.000 131.850 169.410 ;
        RECT 132.190 168.540 132.360 168.870 ;
        RECT 132.530 168.840 133.570 169.010 ;
        RECT 132.530 168.400 133.570 168.570 ;
        RECT 133.740 168.540 133.910 168.870 ;
        RECT 134.250 168.000 134.420 169.410 ;
        RECT 131.550 167.860 134.420 168.000 ;
        RECT 131.680 167.830 134.420 167.860 ;
        RECT 134.980 169.540 137.810 169.590 ;
        RECT 134.980 169.420 137.930 169.540 ;
        RECT 153.730 169.520 156.470 169.590 ;
        RECT 134.980 168.010 135.150 169.420 ;
        RECT 135.490 168.550 135.660 168.880 ;
        RECT 135.875 168.850 136.915 169.020 ;
        RECT 135.875 168.410 136.915 168.580 ;
        RECT 137.130 168.550 137.300 168.880 ;
        RECT 137.640 168.010 137.930 169.420 ;
        RECT 134.980 167.890 137.930 168.010 ;
        RECT 153.600 169.420 156.470 169.520 ;
        RECT 153.600 168.010 153.900 169.420 ;
        RECT 154.240 168.550 154.410 168.880 ;
        RECT 154.580 168.850 155.620 169.020 ;
        RECT 154.580 168.410 155.620 168.580 ;
        RECT 155.790 168.550 155.960 168.880 ;
        RECT 156.300 168.010 156.470 169.420 ;
        RECT 134.980 167.840 137.810 167.890 ;
        RECT 153.600 167.870 156.470 168.010 ;
        RECT 153.730 167.840 156.470 167.870 ;
        RECT 157.030 169.550 159.860 169.600 ;
        RECT 157.030 169.430 159.980 169.550 ;
        RECT 157.030 168.020 157.200 169.430 ;
        RECT 157.540 168.560 157.710 168.890 ;
        RECT 157.925 168.860 158.965 169.030 ;
        RECT 157.925 168.420 158.965 168.590 ;
        RECT 159.180 168.560 159.350 168.890 ;
        RECT 159.690 168.020 159.980 169.430 ;
        RECT 157.030 167.900 159.980 168.020 ;
        RECT 157.030 167.850 159.860 167.900 ;
        RECT 131.680 167.410 134.420 167.480 ;
        RECT 131.550 167.310 134.420 167.410 ;
        RECT 131.550 165.900 131.850 167.310 ;
        RECT 132.190 166.440 132.360 166.770 ;
        RECT 132.530 166.740 133.570 166.910 ;
        RECT 132.530 166.300 133.570 166.470 ;
        RECT 133.740 166.440 133.910 166.770 ;
        RECT 134.250 165.900 134.420 167.310 ;
        RECT 131.550 165.760 134.420 165.900 ;
        RECT 131.680 165.730 134.420 165.760 ;
        RECT 134.980 167.440 137.810 167.490 ;
        RECT 134.980 167.320 137.930 167.440 ;
        RECT 153.730 167.420 156.470 167.490 ;
        RECT 134.980 165.910 135.150 167.320 ;
        RECT 135.490 166.450 135.660 166.780 ;
        RECT 135.875 166.750 136.915 166.920 ;
        RECT 135.875 166.310 136.915 166.480 ;
        RECT 137.130 166.450 137.300 166.780 ;
        RECT 137.640 165.910 137.930 167.320 ;
        RECT 134.980 165.790 137.930 165.910 ;
        RECT 153.600 167.320 156.470 167.420 ;
        RECT 153.600 165.910 153.900 167.320 ;
        RECT 154.240 166.450 154.410 166.780 ;
        RECT 154.580 166.750 155.620 166.920 ;
        RECT 154.580 166.310 155.620 166.480 ;
        RECT 155.790 166.450 155.960 166.780 ;
        RECT 156.300 165.910 156.470 167.320 ;
        RECT 134.980 165.740 137.810 165.790 ;
        RECT 153.600 165.770 156.470 165.910 ;
        RECT 153.730 165.740 156.470 165.770 ;
        RECT 157.030 167.450 159.860 167.500 ;
        RECT 157.030 167.330 159.980 167.450 ;
        RECT 157.030 165.920 157.200 167.330 ;
        RECT 157.540 166.460 157.710 166.790 ;
        RECT 157.925 166.760 158.965 166.930 ;
        RECT 157.925 166.320 158.965 166.490 ;
        RECT 159.180 166.460 159.350 166.790 ;
        RECT 159.690 165.920 159.980 167.330 ;
        RECT 157.030 165.800 159.980 165.920 ;
        RECT 157.030 165.750 159.860 165.800 ;
        RECT 131.680 165.310 134.420 165.380 ;
        RECT 131.550 165.210 134.420 165.310 ;
        RECT 131.550 163.800 131.850 165.210 ;
        RECT 132.190 164.340 132.360 164.670 ;
        RECT 132.530 164.640 133.570 164.810 ;
        RECT 132.530 164.200 133.570 164.370 ;
        RECT 133.740 164.340 133.910 164.670 ;
        RECT 134.250 163.800 134.420 165.210 ;
        RECT 131.550 163.660 134.420 163.800 ;
        RECT 131.680 163.630 134.420 163.660 ;
        RECT 134.980 165.340 137.810 165.390 ;
        RECT 134.980 165.220 137.930 165.340 ;
        RECT 153.730 165.320 156.470 165.390 ;
        RECT 134.980 163.810 135.150 165.220 ;
        RECT 135.490 164.350 135.660 164.680 ;
        RECT 135.875 164.650 136.915 164.820 ;
        RECT 135.875 164.210 136.915 164.380 ;
        RECT 137.130 164.350 137.300 164.680 ;
        RECT 137.640 163.810 137.930 165.220 ;
        RECT 134.980 163.690 137.930 163.810 ;
        RECT 153.600 165.220 156.470 165.320 ;
        RECT 153.600 163.810 153.900 165.220 ;
        RECT 154.240 164.350 154.410 164.680 ;
        RECT 154.580 164.650 155.620 164.820 ;
        RECT 154.580 164.210 155.620 164.380 ;
        RECT 155.790 164.350 155.960 164.680 ;
        RECT 156.300 163.810 156.470 165.220 ;
        RECT 134.980 163.640 137.810 163.690 ;
        RECT 153.600 163.670 156.470 163.810 ;
        RECT 153.730 163.640 156.470 163.670 ;
        RECT 157.030 165.350 159.860 165.400 ;
        RECT 157.030 165.230 159.980 165.350 ;
        RECT 157.030 163.820 157.200 165.230 ;
        RECT 157.540 164.360 157.710 164.690 ;
        RECT 157.925 164.660 158.965 164.830 ;
        RECT 157.925 164.220 158.965 164.390 ;
        RECT 159.180 164.360 159.350 164.690 ;
        RECT 159.690 163.820 159.980 165.230 ;
        RECT 157.030 163.700 159.980 163.820 ;
        RECT 157.030 163.650 159.860 163.700 ;
        RECT 131.680 163.210 134.420 163.280 ;
        RECT 131.550 163.110 134.420 163.210 ;
        RECT 131.550 161.700 131.850 163.110 ;
        RECT 132.190 162.240 132.360 162.570 ;
        RECT 132.530 162.540 133.570 162.710 ;
        RECT 132.530 162.100 133.570 162.270 ;
        RECT 133.740 162.240 133.910 162.570 ;
        RECT 134.250 161.700 134.420 163.110 ;
        RECT 131.550 161.560 134.420 161.700 ;
        RECT 131.680 161.530 134.420 161.560 ;
        RECT 134.980 163.240 137.810 163.290 ;
        RECT 134.980 163.120 137.930 163.240 ;
        RECT 153.730 163.220 156.470 163.290 ;
        RECT 134.980 161.710 135.150 163.120 ;
        RECT 135.490 162.250 135.660 162.580 ;
        RECT 135.875 162.550 136.915 162.720 ;
        RECT 135.875 162.110 136.915 162.280 ;
        RECT 137.130 162.250 137.300 162.580 ;
        RECT 137.640 161.710 137.930 163.120 ;
        RECT 134.980 161.590 137.930 161.710 ;
        RECT 153.600 163.120 156.470 163.220 ;
        RECT 153.600 161.710 153.900 163.120 ;
        RECT 154.240 162.250 154.410 162.580 ;
        RECT 154.580 162.550 155.620 162.720 ;
        RECT 154.580 162.110 155.620 162.280 ;
        RECT 155.790 162.250 155.960 162.580 ;
        RECT 156.300 161.710 156.470 163.120 ;
        RECT 134.980 161.540 137.810 161.590 ;
        RECT 153.600 161.570 156.470 161.710 ;
        RECT 153.730 161.540 156.470 161.570 ;
        RECT 157.030 163.250 159.860 163.300 ;
        RECT 157.030 163.130 159.980 163.250 ;
        RECT 157.030 161.720 157.200 163.130 ;
        RECT 157.540 162.260 157.710 162.590 ;
        RECT 157.925 162.560 158.965 162.730 ;
        RECT 157.925 162.120 158.965 162.290 ;
        RECT 159.180 162.260 159.350 162.590 ;
        RECT 159.690 161.720 159.980 163.130 ;
        RECT 157.030 161.600 159.980 161.720 ;
        RECT 157.030 161.550 159.860 161.600 ;
        RECT 131.680 161.110 134.420 161.180 ;
        RECT 131.550 161.010 134.420 161.110 ;
        RECT 131.550 159.600 131.850 161.010 ;
        RECT 132.190 160.140 132.360 160.470 ;
        RECT 132.530 160.440 133.570 160.610 ;
        RECT 132.530 160.000 133.570 160.170 ;
        RECT 133.740 160.140 133.910 160.470 ;
        RECT 134.250 159.600 134.420 161.010 ;
        RECT 131.550 159.460 134.420 159.600 ;
        RECT 131.680 159.430 134.420 159.460 ;
        RECT 134.980 161.140 137.810 161.190 ;
        RECT 134.980 161.020 137.930 161.140 ;
        RECT 153.730 161.120 156.470 161.190 ;
        RECT 134.980 159.610 135.150 161.020 ;
        RECT 135.490 160.150 135.660 160.480 ;
        RECT 135.875 160.450 136.915 160.620 ;
        RECT 135.875 160.010 136.915 160.180 ;
        RECT 137.130 160.150 137.300 160.480 ;
        RECT 137.640 159.610 137.930 161.020 ;
        RECT 134.980 159.490 137.930 159.610 ;
        RECT 153.600 161.020 156.470 161.120 ;
        RECT 153.600 159.610 153.900 161.020 ;
        RECT 154.240 160.150 154.410 160.480 ;
        RECT 154.580 160.450 155.620 160.620 ;
        RECT 154.580 160.010 155.620 160.180 ;
        RECT 155.790 160.150 155.960 160.480 ;
        RECT 156.300 159.610 156.470 161.020 ;
        RECT 134.980 159.440 137.810 159.490 ;
        RECT 153.600 159.470 156.470 159.610 ;
        RECT 153.730 159.440 156.470 159.470 ;
        RECT 157.030 161.150 159.860 161.200 ;
        RECT 157.030 161.030 159.980 161.150 ;
        RECT 157.030 159.620 157.200 161.030 ;
        RECT 157.540 160.160 157.710 160.490 ;
        RECT 157.925 160.460 158.965 160.630 ;
        RECT 157.925 160.020 158.965 160.190 ;
        RECT 159.180 160.160 159.350 160.490 ;
        RECT 159.690 159.620 159.980 161.030 ;
        RECT 157.030 159.500 159.980 159.620 ;
        RECT 157.030 159.450 159.860 159.500 ;
        RECT 131.680 159.010 134.420 159.080 ;
        RECT 131.550 158.910 134.420 159.010 ;
        RECT 131.550 157.500 131.850 158.910 ;
        RECT 132.190 158.040 132.360 158.370 ;
        RECT 132.530 158.340 133.570 158.510 ;
        RECT 132.530 157.900 133.570 158.070 ;
        RECT 133.740 158.040 133.910 158.370 ;
        RECT 134.250 157.500 134.420 158.910 ;
        RECT 131.550 157.360 134.420 157.500 ;
        RECT 131.680 157.330 134.420 157.360 ;
        RECT 134.980 159.040 137.810 159.090 ;
        RECT 134.980 158.920 137.930 159.040 ;
        RECT 153.730 159.020 156.470 159.090 ;
        RECT 134.980 157.510 135.150 158.920 ;
        RECT 135.490 158.050 135.660 158.380 ;
        RECT 135.875 158.350 136.915 158.520 ;
        RECT 135.875 157.910 136.915 158.080 ;
        RECT 137.130 158.050 137.300 158.380 ;
        RECT 137.640 157.510 137.930 158.920 ;
        RECT 134.980 157.390 137.930 157.510 ;
        RECT 153.600 158.920 156.470 159.020 ;
        RECT 153.600 157.510 153.900 158.920 ;
        RECT 154.240 158.050 154.410 158.380 ;
        RECT 154.580 158.350 155.620 158.520 ;
        RECT 154.580 157.910 155.620 158.080 ;
        RECT 155.790 158.050 155.960 158.380 ;
        RECT 156.300 157.510 156.470 158.920 ;
        RECT 134.980 157.340 137.810 157.390 ;
        RECT 153.600 157.370 156.470 157.510 ;
        RECT 153.730 157.340 156.470 157.370 ;
        RECT 157.030 159.050 159.860 159.100 ;
        RECT 157.030 158.930 159.980 159.050 ;
        RECT 157.030 157.520 157.200 158.930 ;
        RECT 157.540 158.060 157.710 158.390 ;
        RECT 157.925 158.360 158.965 158.530 ;
        RECT 157.925 157.920 158.965 158.090 ;
        RECT 159.180 158.060 159.350 158.390 ;
        RECT 159.690 157.520 159.980 158.930 ;
        RECT 157.030 157.400 159.980 157.520 ;
        RECT 157.030 157.350 159.860 157.400 ;
        RECT 131.680 156.910 134.420 156.980 ;
        RECT 131.550 156.810 134.420 156.910 ;
        RECT 131.550 155.400 131.850 156.810 ;
        RECT 132.190 155.940 132.360 156.270 ;
        RECT 132.530 156.240 133.570 156.410 ;
        RECT 132.530 155.800 133.570 155.970 ;
        RECT 133.740 155.940 133.910 156.270 ;
        RECT 134.250 155.400 134.420 156.810 ;
        RECT 131.550 155.260 134.420 155.400 ;
        RECT 131.680 155.230 134.420 155.260 ;
        RECT 134.980 156.940 137.810 156.990 ;
        RECT 134.980 156.820 137.930 156.940 ;
        RECT 153.730 156.920 156.470 156.990 ;
        RECT 134.980 155.410 135.150 156.820 ;
        RECT 135.490 155.950 135.660 156.280 ;
        RECT 135.875 156.250 136.915 156.420 ;
        RECT 135.875 155.810 136.915 155.980 ;
        RECT 137.130 155.950 137.300 156.280 ;
        RECT 137.640 155.410 137.930 156.820 ;
        RECT 134.980 155.290 137.930 155.410 ;
        RECT 153.600 156.820 156.470 156.920 ;
        RECT 153.600 155.410 153.900 156.820 ;
        RECT 154.240 155.950 154.410 156.280 ;
        RECT 154.580 156.250 155.620 156.420 ;
        RECT 154.580 155.810 155.620 155.980 ;
        RECT 155.790 155.950 155.960 156.280 ;
        RECT 156.300 155.410 156.470 156.820 ;
        RECT 134.980 155.240 137.810 155.290 ;
        RECT 153.600 155.270 156.470 155.410 ;
        RECT 153.730 155.240 156.470 155.270 ;
        RECT 157.030 156.950 159.860 157.000 ;
        RECT 157.030 156.830 159.980 156.950 ;
        RECT 157.030 155.420 157.200 156.830 ;
        RECT 157.540 155.960 157.710 156.290 ;
        RECT 157.925 156.260 158.965 156.430 ;
        RECT 157.925 155.820 158.965 155.990 ;
        RECT 159.180 155.960 159.350 156.290 ;
        RECT 159.690 155.420 159.980 156.830 ;
        RECT 157.030 155.300 159.980 155.420 ;
        RECT 157.030 155.250 159.860 155.300 ;
        RECT 131.680 154.810 134.420 154.880 ;
        RECT 131.550 154.710 134.420 154.810 ;
        RECT 131.550 153.300 131.850 154.710 ;
        RECT 132.190 153.840 132.360 154.170 ;
        RECT 132.530 154.140 133.570 154.310 ;
        RECT 132.530 153.700 133.570 153.870 ;
        RECT 133.740 153.840 133.910 154.170 ;
        RECT 134.250 153.300 134.420 154.710 ;
        RECT 131.550 153.160 134.420 153.300 ;
        RECT 131.680 153.130 134.420 153.160 ;
        RECT 134.980 154.840 137.810 154.890 ;
        RECT 134.980 154.720 137.930 154.840 ;
        RECT 153.730 154.820 156.470 154.890 ;
        RECT 134.980 153.310 135.150 154.720 ;
        RECT 135.490 153.850 135.660 154.180 ;
        RECT 135.875 154.150 136.915 154.320 ;
        RECT 135.875 153.710 136.915 153.880 ;
        RECT 137.130 153.850 137.300 154.180 ;
        RECT 137.640 153.310 137.930 154.720 ;
        RECT 134.980 153.190 137.930 153.310 ;
        RECT 153.600 154.720 156.470 154.820 ;
        RECT 153.600 153.310 153.900 154.720 ;
        RECT 154.240 153.850 154.410 154.180 ;
        RECT 154.580 154.150 155.620 154.320 ;
        RECT 154.580 153.710 155.620 153.880 ;
        RECT 155.790 153.850 155.960 154.180 ;
        RECT 156.300 153.310 156.470 154.720 ;
        RECT 134.980 153.140 137.810 153.190 ;
        RECT 153.600 153.170 156.470 153.310 ;
        RECT 153.730 153.140 156.470 153.170 ;
        RECT 157.030 154.850 159.860 154.900 ;
        RECT 157.030 154.730 159.980 154.850 ;
        RECT 157.030 153.320 157.200 154.730 ;
        RECT 157.540 153.860 157.710 154.190 ;
        RECT 157.925 154.160 158.965 154.330 ;
        RECT 157.925 153.720 158.965 153.890 ;
        RECT 159.180 153.860 159.350 154.190 ;
        RECT 159.690 153.320 159.980 154.730 ;
        RECT 157.030 153.200 159.980 153.320 ;
        RECT 157.030 153.150 159.860 153.200 ;
        RECT 131.680 152.710 134.420 152.780 ;
        RECT 131.550 152.610 134.420 152.710 ;
        RECT 131.550 151.200 131.850 152.610 ;
        RECT 132.190 151.740 132.360 152.070 ;
        RECT 132.530 152.040 133.570 152.210 ;
        RECT 132.530 151.600 133.570 151.770 ;
        RECT 133.740 151.740 133.910 152.070 ;
        RECT 134.250 151.200 134.420 152.610 ;
        RECT 131.550 151.060 134.420 151.200 ;
        RECT 131.680 151.030 134.420 151.060 ;
        RECT 134.980 152.740 137.810 152.790 ;
        RECT 134.980 152.620 137.930 152.740 ;
        RECT 153.730 152.720 156.470 152.790 ;
        RECT 134.980 151.210 135.150 152.620 ;
        RECT 135.490 151.750 135.660 152.080 ;
        RECT 135.875 152.050 136.915 152.220 ;
        RECT 135.875 151.610 136.915 151.780 ;
        RECT 137.130 151.750 137.300 152.080 ;
        RECT 137.640 151.210 137.930 152.620 ;
        RECT 134.980 151.090 137.930 151.210 ;
        RECT 153.600 152.620 156.470 152.720 ;
        RECT 153.600 151.210 153.900 152.620 ;
        RECT 154.240 151.750 154.410 152.080 ;
        RECT 154.580 152.050 155.620 152.220 ;
        RECT 154.580 151.610 155.620 151.780 ;
        RECT 155.790 151.750 155.960 152.080 ;
        RECT 156.300 151.210 156.470 152.620 ;
        RECT 134.980 151.040 137.810 151.090 ;
        RECT 153.600 151.070 156.470 151.210 ;
        RECT 153.730 151.040 156.470 151.070 ;
        RECT 157.030 152.750 159.860 152.800 ;
        RECT 157.030 152.630 159.980 152.750 ;
        RECT 157.030 151.220 157.200 152.630 ;
        RECT 157.540 151.760 157.710 152.090 ;
        RECT 157.925 152.060 158.965 152.230 ;
        RECT 157.925 151.620 158.965 151.790 ;
        RECT 159.180 151.760 159.350 152.090 ;
        RECT 159.690 151.220 159.980 152.630 ;
        RECT 157.030 151.100 159.980 151.220 ;
        RECT 157.030 151.050 159.860 151.100 ;
        RECT 131.680 150.610 134.420 150.680 ;
        RECT 131.550 150.510 134.420 150.610 ;
        RECT 131.550 149.100 131.850 150.510 ;
        RECT 132.190 149.640 132.360 149.970 ;
        RECT 132.530 149.940 133.570 150.110 ;
        RECT 132.530 149.500 133.570 149.670 ;
        RECT 133.740 149.640 133.910 149.970 ;
        RECT 134.250 149.100 134.420 150.510 ;
        RECT 131.550 148.960 134.420 149.100 ;
        RECT 131.680 148.930 134.420 148.960 ;
        RECT 134.980 150.640 137.810 150.690 ;
        RECT 134.980 150.520 137.930 150.640 ;
        RECT 153.730 150.620 156.470 150.690 ;
        RECT 134.980 149.110 135.150 150.520 ;
        RECT 135.490 149.650 135.660 149.980 ;
        RECT 135.875 149.950 136.915 150.120 ;
        RECT 135.875 149.510 136.915 149.680 ;
        RECT 137.130 149.650 137.300 149.980 ;
        RECT 137.640 149.110 137.930 150.520 ;
        RECT 134.980 148.990 137.930 149.110 ;
        RECT 153.600 150.520 156.470 150.620 ;
        RECT 153.600 149.110 153.900 150.520 ;
        RECT 154.240 149.650 154.410 149.980 ;
        RECT 154.580 149.950 155.620 150.120 ;
        RECT 154.580 149.510 155.620 149.680 ;
        RECT 155.790 149.650 155.960 149.980 ;
        RECT 156.300 149.110 156.470 150.520 ;
        RECT 134.980 148.940 137.810 148.990 ;
        RECT 153.600 148.970 156.470 149.110 ;
        RECT 153.730 148.940 156.470 148.970 ;
        RECT 157.030 150.650 159.860 150.700 ;
        RECT 157.030 150.530 159.980 150.650 ;
        RECT 157.030 149.120 157.200 150.530 ;
        RECT 157.540 149.660 157.710 149.990 ;
        RECT 157.925 149.960 158.965 150.130 ;
        RECT 157.925 149.520 158.965 149.690 ;
        RECT 159.180 149.660 159.350 149.990 ;
        RECT 159.690 149.120 159.980 150.530 ;
        RECT 157.030 149.000 159.980 149.120 ;
        RECT 157.030 148.950 159.860 149.000 ;
        RECT 131.680 148.510 134.420 148.580 ;
        RECT 131.550 148.410 134.420 148.510 ;
        RECT 131.550 147.000 131.850 148.410 ;
        RECT 132.190 147.540 132.360 147.870 ;
        RECT 132.530 147.840 133.570 148.010 ;
        RECT 132.530 147.400 133.570 147.570 ;
        RECT 133.740 147.540 133.910 147.870 ;
        RECT 134.250 147.000 134.420 148.410 ;
        RECT 131.550 146.860 134.420 147.000 ;
        RECT 131.680 146.830 134.420 146.860 ;
        RECT 134.980 148.540 137.810 148.590 ;
        RECT 134.980 148.420 137.930 148.540 ;
        RECT 153.730 148.520 156.470 148.590 ;
        RECT 134.980 147.010 135.150 148.420 ;
        RECT 135.490 147.550 135.660 147.880 ;
        RECT 135.875 147.850 136.915 148.020 ;
        RECT 135.875 147.410 136.915 147.580 ;
        RECT 137.130 147.550 137.300 147.880 ;
        RECT 137.640 147.010 137.930 148.420 ;
        RECT 134.980 146.890 137.930 147.010 ;
        RECT 153.600 148.420 156.470 148.520 ;
        RECT 153.600 147.010 153.900 148.420 ;
        RECT 154.240 147.550 154.410 147.880 ;
        RECT 154.580 147.850 155.620 148.020 ;
        RECT 154.580 147.410 155.620 147.580 ;
        RECT 155.790 147.550 155.960 147.880 ;
        RECT 156.300 147.010 156.470 148.420 ;
        RECT 134.980 146.840 137.810 146.890 ;
        RECT 153.600 146.870 156.470 147.010 ;
        RECT 153.730 146.840 156.470 146.870 ;
        RECT 157.030 148.550 159.860 148.600 ;
        RECT 157.030 148.430 159.980 148.550 ;
        RECT 157.030 147.020 157.200 148.430 ;
        RECT 157.540 147.560 157.710 147.890 ;
        RECT 157.925 147.860 158.965 148.030 ;
        RECT 157.925 147.420 158.965 147.590 ;
        RECT 159.180 147.560 159.350 147.890 ;
        RECT 159.690 147.020 159.980 148.430 ;
        RECT 157.030 146.900 159.980 147.020 ;
        RECT 157.030 146.850 159.860 146.900 ;
        RECT 131.680 146.410 134.420 146.480 ;
        RECT 131.550 146.310 134.420 146.410 ;
        RECT 131.550 144.900 131.850 146.310 ;
        RECT 132.190 145.440 132.360 145.770 ;
        RECT 132.530 145.740 133.570 145.910 ;
        RECT 132.530 145.300 133.570 145.470 ;
        RECT 133.740 145.440 133.910 145.770 ;
        RECT 134.250 144.900 134.420 146.310 ;
        RECT 131.550 144.760 134.420 144.900 ;
        RECT 131.680 144.730 134.420 144.760 ;
        RECT 134.980 146.440 137.810 146.490 ;
        RECT 134.980 146.320 137.930 146.440 ;
        RECT 153.730 146.420 156.470 146.490 ;
        RECT 134.980 144.910 135.150 146.320 ;
        RECT 135.490 145.450 135.660 145.780 ;
        RECT 135.875 145.750 136.915 145.920 ;
        RECT 135.875 145.310 136.915 145.480 ;
        RECT 137.130 145.450 137.300 145.780 ;
        RECT 137.640 144.910 137.930 146.320 ;
        RECT 134.980 144.790 137.930 144.910 ;
        RECT 153.600 146.320 156.470 146.420 ;
        RECT 153.600 144.910 153.900 146.320 ;
        RECT 154.240 145.450 154.410 145.780 ;
        RECT 154.580 145.750 155.620 145.920 ;
        RECT 154.580 145.310 155.620 145.480 ;
        RECT 155.790 145.450 155.960 145.780 ;
        RECT 156.300 144.910 156.470 146.320 ;
        RECT 134.980 144.740 137.810 144.790 ;
        RECT 153.600 144.770 156.470 144.910 ;
        RECT 153.730 144.740 156.470 144.770 ;
        RECT 157.030 146.450 159.860 146.500 ;
        RECT 157.030 146.330 159.980 146.450 ;
        RECT 157.030 144.920 157.200 146.330 ;
        RECT 157.540 145.460 157.710 145.790 ;
        RECT 157.925 145.760 158.965 145.930 ;
        RECT 157.925 145.320 158.965 145.490 ;
        RECT 159.180 145.460 159.350 145.790 ;
        RECT 159.690 144.920 159.980 146.330 ;
        RECT 157.030 144.800 159.980 144.920 ;
        RECT 157.030 144.750 159.860 144.800 ;
        RECT 131.680 144.310 134.420 144.380 ;
        RECT 131.550 144.210 134.420 144.310 ;
        RECT 131.550 142.800 131.850 144.210 ;
        RECT 132.190 143.340 132.360 143.670 ;
        RECT 132.530 143.640 133.570 143.810 ;
        RECT 132.530 143.200 133.570 143.370 ;
        RECT 133.740 143.340 133.910 143.670 ;
        RECT 134.250 142.800 134.420 144.210 ;
        RECT 131.550 142.660 134.420 142.800 ;
        RECT 131.680 142.630 134.420 142.660 ;
        RECT 134.980 144.340 137.810 144.390 ;
        RECT 134.980 144.220 137.930 144.340 ;
        RECT 153.730 144.320 156.470 144.390 ;
        RECT 134.980 142.810 135.150 144.220 ;
        RECT 135.490 143.350 135.660 143.680 ;
        RECT 135.875 143.650 136.915 143.820 ;
        RECT 135.875 143.210 136.915 143.380 ;
        RECT 137.130 143.350 137.300 143.680 ;
        RECT 137.640 142.810 137.930 144.220 ;
        RECT 134.980 142.690 137.930 142.810 ;
        RECT 153.600 144.220 156.470 144.320 ;
        RECT 153.600 142.810 153.900 144.220 ;
        RECT 154.240 143.350 154.410 143.680 ;
        RECT 154.580 143.650 155.620 143.820 ;
        RECT 154.580 143.210 155.620 143.380 ;
        RECT 155.790 143.350 155.960 143.680 ;
        RECT 156.300 142.810 156.470 144.220 ;
        RECT 134.980 142.640 137.810 142.690 ;
        RECT 153.600 142.670 156.470 142.810 ;
        RECT 153.730 142.640 156.470 142.670 ;
        RECT 157.030 144.350 159.860 144.400 ;
        RECT 157.030 144.230 159.980 144.350 ;
        RECT 157.030 142.820 157.200 144.230 ;
        RECT 157.540 143.360 157.710 143.690 ;
        RECT 157.925 143.660 158.965 143.830 ;
        RECT 157.925 143.220 158.965 143.390 ;
        RECT 159.180 143.360 159.350 143.690 ;
        RECT 159.690 142.820 159.980 144.230 ;
        RECT 157.030 142.700 159.980 142.820 ;
        RECT 157.030 142.650 159.860 142.700 ;
        RECT 131.680 142.210 134.420 142.280 ;
        RECT 131.550 142.110 134.420 142.210 ;
        RECT 131.550 140.700 131.850 142.110 ;
        RECT 132.190 141.240 132.360 141.570 ;
        RECT 132.530 141.540 133.570 141.710 ;
        RECT 132.530 141.100 133.570 141.270 ;
        RECT 133.740 141.240 133.910 141.570 ;
        RECT 134.250 140.700 134.420 142.110 ;
        RECT 131.550 140.560 134.420 140.700 ;
        RECT 131.680 140.530 134.420 140.560 ;
        RECT 134.980 142.240 137.810 142.290 ;
        RECT 134.980 142.120 137.930 142.240 ;
        RECT 153.730 142.220 156.470 142.290 ;
        RECT 134.980 140.710 135.150 142.120 ;
        RECT 135.490 141.250 135.660 141.580 ;
        RECT 135.875 141.550 136.915 141.720 ;
        RECT 135.875 141.110 136.915 141.280 ;
        RECT 137.130 141.250 137.300 141.580 ;
        RECT 137.640 140.710 137.930 142.120 ;
        RECT 134.980 140.590 137.930 140.710 ;
        RECT 153.600 142.120 156.470 142.220 ;
        RECT 153.600 140.710 153.900 142.120 ;
        RECT 154.240 141.250 154.410 141.580 ;
        RECT 154.580 141.550 155.620 141.720 ;
        RECT 154.580 141.110 155.620 141.280 ;
        RECT 155.790 141.250 155.960 141.580 ;
        RECT 156.300 140.710 156.470 142.120 ;
        RECT 134.980 140.540 137.810 140.590 ;
        RECT 153.600 140.570 156.470 140.710 ;
        RECT 153.730 140.540 156.470 140.570 ;
        RECT 157.030 142.250 159.860 142.300 ;
        RECT 157.030 142.130 159.980 142.250 ;
        RECT 157.030 140.720 157.200 142.130 ;
        RECT 157.540 141.260 157.710 141.590 ;
        RECT 157.925 141.560 158.965 141.730 ;
        RECT 157.925 141.120 158.965 141.290 ;
        RECT 159.180 141.260 159.350 141.590 ;
        RECT 159.690 140.720 159.980 142.130 ;
        RECT 157.030 140.600 159.980 140.720 ;
        RECT 157.030 140.550 159.860 140.600 ;
        RECT 131.680 140.110 134.420 140.180 ;
        RECT 131.550 140.010 134.420 140.110 ;
        RECT 131.550 138.600 131.850 140.010 ;
        RECT 132.190 139.140 132.360 139.470 ;
        RECT 132.530 139.440 133.570 139.610 ;
        RECT 132.530 139.000 133.570 139.170 ;
        RECT 133.740 139.140 133.910 139.470 ;
        RECT 134.250 138.600 134.420 140.010 ;
        RECT 131.550 138.460 134.420 138.600 ;
        RECT 131.680 138.430 134.420 138.460 ;
        RECT 134.980 140.140 137.810 140.190 ;
        RECT 134.980 140.020 137.930 140.140 ;
        RECT 153.730 140.120 156.470 140.190 ;
        RECT 134.980 138.610 135.150 140.020 ;
        RECT 135.490 139.150 135.660 139.480 ;
        RECT 135.875 139.450 136.915 139.620 ;
        RECT 135.875 139.010 136.915 139.180 ;
        RECT 137.130 139.150 137.300 139.480 ;
        RECT 137.640 138.610 137.930 140.020 ;
        RECT 134.980 138.490 137.930 138.610 ;
        RECT 153.600 140.020 156.470 140.120 ;
        RECT 153.600 138.610 153.900 140.020 ;
        RECT 154.240 139.150 154.410 139.480 ;
        RECT 154.580 139.450 155.620 139.620 ;
        RECT 154.580 139.010 155.620 139.180 ;
        RECT 155.790 139.150 155.960 139.480 ;
        RECT 156.300 138.610 156.470 140.020 ;
        RECT 134.980 138.440 137.810 138.490 ;
        RECT 153.600 138.470 156.470 138.610 ;
        RECT 153.730 138.440 156.470 138.470 ;
        RECT 157.030 140.150 159.860 140.200 ;
        RECT 157.030 140.030 159.980 140.150 ;
        RECT 157.030 138.620 157.200 140.030 ;
        RECT 157.540 139.160 157.710 139.490 ;
        RECT 157.925 139.460 158.965 139.630 ;
        RECT 157.925 139.020 158.965 139.190 ;
        RECT 159.180 139.160 159.350 139.490 ;
        RECT 159.690 138.620 159.980 140.030 ;
        RECT 157.030 138.500 159.980 138.620 ;
        RECT 157.030 138.450 159.860 138.500 ;
        RECT 131.680 138.010 134.420 138.080 ;
        RECT 131.550 137.910 134.420 138.010 ;
        RECT 131.550 136.500 131.850 137.910 ;
        RECT 132.190 137.040 132.360 137.370 ;
        RECT 132.530 137.340 133.570 137.510 ;
        RECT 132.530 136.900 133.570 137.070 ;
        RECT 133.740 137.040 133.910 137.370 ;
        RECT 134.250 136.500 134.420 137.910 ;
        RECT 131.550 136.360 134.420 136.500 ;
        RECT 131.680 136.330 134.420 136.360 ;
        RECT 134.980 138.040 137.810 138.090 ;
        RECT 134.980 137.920 137.930 138.040 ;
        RECT 153.730 138.020 156.470 138.090 ;
        RECT 134.980 136.510 135.150 137.920 ;
        RECT 135.490 137.050 135.660 137.380 ;
        RECT 135.875 137.350 136.915 137.520 ;
        RECT 135.875 136.910 136.915 137.080 ;
        RECT 137.130 137.050 137.300 137.380 ;
        RECT 137.640 136.510 137.930 137.920 ;
        RECT 134.980 136.390 137.930 136.510 ;
        RECT 153.600 137.920 156.470 138.020 ;
        RECT 153.600 136.510 153.900 137.920 ;
        RECT 154.240 137.050 154.410 137.380 ;
        RECT 154.580 137.350 155.620 137.520 ;
        RECT 154.580 136.910 155.620 137.080 ;
        RECT 155.790 137.050 155.960 137.380 ;
        RECT 156.300 136.510 156.470 137.920 ;
        RECT 134.980 136.340 137.810 136.390 ;
        RECT 153.600 136.370 156.470 136.510 ;
        RECT 153.730 136.340 156.470 136.370 ;
        RECT 157.030 138.050 159.860 138.100 ;
        RECT 157.030 137.930 159.980 138.050 ;
        RECT 157.030 136.520 157.200 137.930 ;
        RECT 157.540 137.060 157.710 137.390 ;
        RECT 157.925 137.360 158.965 137.530 ;
        RECT 157.925 136.920 158.965 137.090 ;
        RECT 159.180 137.060 159.350 137.390 ;
        RECT 159.690 136.520 159.980 137.930 ;
        RECT 157.030 136.400 159.980 136.520 ;
        RECT 157.030 136.350 159.860 136.400 ;
        RECT 131.680 135.910 134.420 135.980 ;
        RECT 131.550 135.810 134.420 135.910 ;
        RECT 131.550 134.400 131.850 135.810 ;
        RECT 132.190 134.940 132.360 135.270 ;
        RECT 132.530 135.240 133.570 135.410 ;
        RECT 132.530 134.800 133.570 134.970 ;
        RECT 133.740 134.940 133.910 135.270 ;
        RECT 134.250 134.400 134.420 135.810 ;
        RECT 131.550 134.260 134.420 134.400 ;
        RECT 131.680 134.230 134.420 134.260 ;
        RECT 134.980 135.940 137.810 135.990 ;
        RECT 134.980 135.820 137.930 135.940 ;
        RECT 153.730 135.920 156.470 135.990 ;
        RECT 134.980 134.410 135.150 135.820 ;
        RECT 135.490 134.950 135.660 135.280 ;
        RECT 135.875 135.250 136.915 135.420 ;
        RECT 135.875 134.810 136.915 134.980 ;
        RECT 137.130 134.950 137.300 135.280 ;
        RECT 137.640 134.410 137.930 135.820 ;
        RECT 134.980 134.290 137.930 134.410 ;
        RECT 153.600 135.820 156.470 135.920 ;
        RECT 153.600 134.410 153.900 135.820 ;
        RECT 154.240 134.950 154.410 135.280 ;
        RECT 154.580 135.250 155.620 135.420 ;
        RECT 154.580 134.810 155.620 134.980 ;
        RECT 155.790 134.950 155.960 135.280 ;
        RECT 156.300 134.410 156.470 135.820 ;
        RECT 134.980 134.240 137.810 134.290 ;
        RECT 153.600 134.270 156.470 134.410 ;
        RECT 153.730 134.240 156.470 134.270 ;
        RECT 157.030 135.950 159.860 136.000 ;
        RECT 157.030 135.830 159.980 135.950 ;
        RECT 157.030 134.420 157.200 135.830 ;
        RECT 157.540 134.960 157.710 135.290 ;
        RECT 157.925 135.260 158.965 135.430 ;
        RECT 157.925 134.820 158.965 134.990 ;
        RECT 159.180 134.960 159.350 135.290 ;
        RECT 159.690 134.420 159.980 135.830 ;
        RECT 157.030 134.300 159.980 134.420 ;
        RECT 157.030 134.250 159.860 134.300 ;
        RECT 131.680 133.810 134.420 133.880 ;
        RECT 131.550 133.710 134.420 133.810 ;
        RECT 131.550 132.300 131.850 133.710 ;
        RECT 132.190 132.840 132.360 133.170 ;
        RECT 132.530 133.140 133.570 133.310 ;
        RECT 132.530 132.700 133.570 132.870 ;
        RECT 133.740 132.840 133.910 133.170 ;
        RECT 134.250 132.300 134.420 133.710 ;
        RECT 131.550 132.160 134.420 132.300 ;
        RECT 131.680 132.130 134.420 132.160 ;
        RECT 134.980 133.840 137.810 133.890 ;
        RECT 134.980 133.720 137.930 133.840 ;
        RECT 153.730 133.820 156.470 133.890 ;
        RECT 134.980 132.310 135.150 133.720 ;
        RECT 135.490 132.850 135.660 133.180 ;
        RECT 135.875 133.150 136.915 133.320 ;
        RECT 135.875 132.710 136.915 132.880 ;
        RECT 137.130 132.850 137.300 133.180 ;
        RECT 137.640 132.310 137.930 133.720 ;
        RECT 134.980 132.190 137.930 132.310 ;
        RECT 153.600 133.720 156.470 133.820 ;
        RECT 153.600 132.310 153.900 133.720 ;
        RECT 154.240 132.850 154.410 133.180 ;
        RECT 154.580 133.150 155.620 133.320 ;
        RECT 154.580 132.710 155.620 132.880 ;
        RECT 155.790 132.850 155.960 133.180 ;
        RECT 156.300 132.310 156.470 133.720 ;
        RECT 134.980 132.140 137.810 132.190 ;
        RECT 153.600 132.170 156.470 132.310 ;
        RECT 153.730 132.140 156.470 132.170 ;
        RECT 157.030 133.850 159.860 133.900 ;
        RECT 157.030 133.730 159.980 133.850 ;
        RECT 157.030 132.320 157.200 133.730 ;
        RECT 157.540 132.860 157.710 133.190 ;
        RECT 157.925 133.160 158.965 133.330 ;
        RECT 157.925 132.720 158.965 132.890 ;
        RECT 159.180 132.860 159.350 133.190 ;
        RECT 159.690 132.320 159.980 133.730 ;
        RECT 157.030 132.200 159.980 132.320 ;
        RECT 157.030 132.150 159.860 132.200 ;
        RECT 131.680 131.710 134.420 131.780 ;
        RECT 131.550 131.610 134.420 131.710 ;
        RECT 131.550 130.200 131.850 131.610 ;
        RECT 132.190 130.740 132.360 131.070 ;
        RECT 132.530 131.040 133.570 131.210 ;
        RECT 132.530 130.600 133.570 130.770 ;
        RECT 133.740 130.740 133.910 131.070 ;
        RECT 134.250 130.200 134.420 131.610 ;
        RECT 131.550 130.060 134.420 130.200 ;
        RECT 131.680 130.030 134.420 130.060 ;
        RECT 134.980 131.740 137.810 131.790 ;
        RECT 134.980 131.620 137.930 131.740 ;
        RECT 153.730 131.720 156.470 131.790 ;
        RECT 134.980 130.210 135.150 131.620 ;
        RECT 135.490 130.750 135.660 131.080 ;
        RECT 135.875 131.050 136.915 131.220 ;
        RECT 135.875 130.610 136.915 130.780 ;
        RECT 137.130 130.750 137.300 131.080 ;
        RECT 137.640 130.210 137.930 131.620 ;
        RECT 134.980 130.090 137.930 130.210 ;
        RECT 153.600 131.620 156.470 131.720 ;
        RECT 153.600 130.210 153.900 131.620 ;
        RECT 154.240 130.750 154.410 131.080 ;
        RECT 154.580 131.050 155.620 131.220 ;
        RECT 154.580 130.610 155.620 130.780 ;
        RECT 155.790 130.750 155.960 131.080 ;
        RECT 156.300 130.210 156.470 131.620 ;
        RECT 134.980 130.040 137.810 130.090 ;
        RECT 153.600 130.070 156.470 130.210 ;
        RECT 153.730 130.040 156.470 130.070 ;
        RECT 157.030 131.750 159.860 131.800 ;
        RECT 157.030 131.630 159.980 131.750 ;
        RECT 157.030 130.220 157.200 131.630 ;
        RECT 157.540 130.760 157.710 131.090 ;
        RECT 157.925 131.060 158.965 131.230 ;
        RECT 157.925 130.620 158.965 130.790 ;
        RECT 159.180 130.760 159.350 131.090 ;
        RECT 159.690 130.220 159.980 131.630 ;
        RECT 157.030 130.100 159.980 130.220 ;
        RECT 157.030 130.050 159.860 130.100 ;
        RECT 131.680 129.610 134.420 129.680 ;
        RECT 131.550 129.510 134.420 129.610 ;
        RECT 131.550 128.100 131.850 129.510 ;
        RECT 132.190 128.640 132.360 128.970 ;
        RECT 132.530 128.940 133.570 129.110 ;
        RECT 132.530 128.500 133.570 128.670 ;
        RECT 133.740 128.640 133.910 128.970 ;
        RECT 134.250 128.100 134.420 129.510 ;
        RECT 131.550 127.960 134.420 128.100 ;
        RECT 131.680 127.930 134.420 127.960 ;
        RECT 134.980 129.640 137.810 129.690 ;
        RECT 134.980 129.520 137.930 129.640 ;
        RECT 153.730 129.620 156.470 129.690 ;
        RECT 134.980 128.110 135.150 129.520 ;
        RECT 135.490 128.650 135.660 128.980 ;
        RECT 135.875 128.950 136.915 129.120 ;
        RECT 135.875 128.510 136.915 128.680 ;
        RECT 137.130 128.650 137.300 128.980 ;
        RECT 137.640 128.110 137.930 129.520 ;
        RECT 134.980 127.990 137.930 128.110 ;
        RECT 153.600 129.520 156.470 129.620 ;
        RECT 153.600 128.110 153.900 129.520 ;
        RECT 154.240 128.650 154.410 128.980 ;
        RECT 154.580 128.950 155.620 129.120 ;
        RECT 154.580 128.510 155.620 128.680 ;
        RECT 155.790 128.650 155.960 128.980 ;
        RECT 156.300 128.110 156.470 129.520 ;
        RECT 134.980 127.940 137.810 127.990 ;
        RECT 153.600 127.970 156.470 128.110 ;
        RECT 153.730 127.940 156.470 127.970 ;
        RECT 157.030 129.650 159.860 129.700 ;
        RECT 157.030 129.530 159.980 129.650 ;
        RECT 157.030 128.120 157.200 129.530 ;
        RECT 157.540 128.660 157.710 128.990 ;
        RECT 157.925 128.960 158.965 129.130 ;
        RECT 157.925 128.520 158.965 128.690 ;
        RECT 159.180 128.660 159.350 128.990 ;
        RECT 159.690 128.120 159.980 129.530 ;
        RECT 157.030 128.000 159.980 128.120 ;
        RECT 157.030 127.950 159.860 128.000 ;
        RECT 131.680 127.510 134.420 127.580 ;
        RECT 131.550 127.410 134.420 127.510 ;
        RECT 131.550 126.000 131.850 127.410 ;
        RECT 132.190 126.540 132.360 126.870 ;
        RECT 132.530 126.840 133.570 127.010 ;
        RECT 132.530 126.400 133.570 126.570 ;
        RECT 133.740 126.540 133.910 126.870 ;
        RECT 134.250 126.000 134.420 127.410 ;
        RECT 131.550 125.860 134.420 126.000 ;
        RECT 131.680 125.830 134.420 125.860 ;
        RECT 134.980 127.540 137.810 127.590 ;
        RECT 134.980 127.420 137.930 127.540 ;
        RECT 153.730 127.520 156.470 127.590 ;
        RECT 134.980 126.010 135.150 127.420 ;
        RECT 135.490 126.550 135.660 126.880 ;
        RECT 135.875 126.850 136.915 127.020 ;
        RECT 135.875 126.410 136.915 126.580 ;
        RECT 137.130 126.550 137.300 126.880 ;
        RECT 137.640 126.010 137.930 127.420 ;
        RECT 134.980 125.890 137.930 126.010 ;
        RECT 153.600 127.420 156.470 127.520 ;
        RECT 153.600 126.010 153.900 127.420 ;
        RECT 154.240 126.550 154.410 126.880 ;
        RECT 154.580 126.850 155.620 127.020 ;
        RECT 154.580 126.410 155.620 126.580 ;
        RECT 155.790 126.550 155.960 126.880 ;
        RECT 156.300 126.010 156.470 127.420 ;
        RECT 134.980 125.840 137.810 125.890 ;
        RECT 153.600 125.870 156.470 126.010 ;
        RECT 153.730 125.840 156.470 125.870 ;
        RECT 157.030 127.550 159.860 127.600 ;
        RECT 157.030 127.430 159.980 127.550 ;
        RECT 157.030 126.020 157.200 127.430 ;
        RECT 157.540 126.560 157.710 126.890 ;
        RECT 157.925 126.860 158.965 127.030 ;
        RECT 157.925 126.420 158.965 126.590 ;
        RECT 159.180 126.560 159.350 126.890 ;
        RECT 159.690 126.020 159.980 127.430 ;
        RECT 157.030 125.900 159.980 126.020 ;
        RECT 157.030 125.850 159.860 125.900 ;
        RECT 131.680 125.410 134.420 125.480 ;
        RECT 131.550 125.310 134.420 125.410 ;
        RECT 131.550 123.900 131.850 125.310 ;
        RECT 132.190 124.440 132.360 124.770 ;
        RECT 132.530 124.740 133.570 124.910 ;
        RECT 132.530 124.300 133.570 124.470 ;
        RECT 133.740 124.440 133.910 124.770 ;
        RECT 134.250 123.900 134.420 125.310 ;
        RECT 131.550 123.760 134.420 123.900 ;
        RECT 131.680 123.730 134.420 123.760 ;
        RECT 134.980 125.440 137.810 125.490 ;
        RECT 134.980 125.320 137.930 125.440 ;
        RECT 153.730 125.420 156.470 125.490 ;
        RECT 134.980 123.910 135.150 125.320 ;
        RECT 135.490 124.450 135.660 124.780 ;
        RECT 135.875 124.750 136.915 124.920 ;
        RECT 135.875 124.310 136.915 124.480 ;
        RECT 137.130 124.450 137.300 124.780 ;
        RECT 137.640 123.910 137.930 125.320 ;
        RECT 134.980 123.790 137.930 123.910 ;
        RECT 153.600 125.320 156.470 125.420 ;
        RECT 153.600 123.910 153.900 125.320 ;
        RECT 154.240 124.450 154.410 124.780 ;
        RECT 154.580 124.750 155.620 124.920 ;
        RECT 154.580 124.310 155.620 124.480 ;
        RECT 155.790 124.450 155.960 124.780 ;
        RECT 156.300 123.910 156.470 125.320 ;
        RECT 134.980 123.740 137.810 123.790 ;
        RECT 153.600 123.770 156.470 123.910 ;
        RECT 153.730 123.740 156.470 123.770 ;
        RECT 157.030 125.450 159.860 125.500 ;
        RECT 157.030 125.330 159.980 125.450 ;
        RECT 157.030 123.920 157.200 125.330 ;
        RECT 157.540 124.460 157.710 124.790 ;
        RECT 157.925 124.760 158.965 124.930 ;
        RECT 157.925 124.320 158.965 124.490 ;
        RECT 159.180 124.460 159.350 124.790 ;
        RECT 159.690 123.920 159.980 125.330 ;
        RECT 157.030 123.800 159.980 123.920 ;
        RECT 157.030 123.750 159.860 123.800 ;
        RECT 131.680 123.310 134.420 123.380 ;
        RECT 131.550 123.210 134.420 123.310 ;
        RECT 131.550 121.800 131.850 123.210 ;
        RECT 132.190 122.340 132.360 122.670 ;
        RECT 132.530 122.640 133.570 122.810 ;
        RECT 132.530 122.200 133.570 122.370 ;
        RECT 133.740 122.340 133.910 122.670 ;
        RECT 134.250 121.800 134.420 123.210 ;
        RECT 131.550 121.660 134.420 121.800 ;
        RECT 131.680 121.630 134.420 121.660 ;
        RECT 134.980 123.340 137.810 123.390 ;
        RECT 134.980 123.220 137.930 123.340 ;
        RECT 153.730 123.320 156.470 123.390 ;
        RECT 134.980 121.810 135.150 123.220 ;
        RECT 135.490 122.350 135.660 122.680 ;
        RECT 135.875 122.650 136.915 122.820 ;
        RECT 135.875 122.210 136.915 122.380 ;
        RECT 137.130 122.350 137.300 122.680 ;
        RECT 137.640 121.810 137.930 123.220 ;
        RECT 134.980 121.690 137.930 121.810 ;
        RECT 153.600 123.220 156.470 123.320 ;
        RECT 153.600 121.810 153.900 123.220 ;
        RECT 154.240 122.350 154.410 122.680 ;
        RECT 154.580 122.650 155.620 122.820 ;
        RECT 154.580 122.210 155.620 122.380 ;
        RECT 155.790 122.350 155.960 122.680 ;
        RECT 156.300 121.810 156.470 123.220 ;
        RECT 134.980 121.640 137.810 121.690 ;
        RECT 153.600 121.670 156.470 121.810 ;
        RECT 153.730 121.640 156.470 121.670 ;
        RECT 157.030 123.350 159.860 123.400 ;
        RECT 157.030 123.230 159.980 123.350 ;
        RECT 157.030 121.820 157.200 123.230 ;
        RECT 157.540 122.360 157.710 122.690 ;
        RECT 157.925 122.660 158.965 122.830 ;
        RECT 157.925 122.220 158.965 122.390 ;
        RECT 159.180 122.360 159.350 122.690 ;
        RECT 159.690 121.820 159.980 123.230 ;
        RECT 157.030 121.700 159.980 121.820 ;
        RECT 157.030 121.650 159.860 121.700 ;
        RECT 131.680 121.210 134.420 121.280 ;
        RECT 131.550 121.110 134.420 121.210 ;
        RECT 131.550 119.700 131.850 121.110 ;
        RECT 132.190 120.240 132.360 120.570 ;
        RECT 132.530 120.540 133.570 120.710 ;
        RECT 132.530 120.100 133.570 120.270 ;
        RECT 133.740 120.240 133.910 120.570 ;
        RECT 134.250 119.700 134.420 121.110 ;
        RECT 131.550 119.560 134.420 119.700 ;
        RECT 131.680 119.530 134.420 119.560 ;
        RECT 134.980 121.240 137.810 121.290 ;
        RECT 134.980 121.120 137.930 121.240 ;
        RECT 153.730 121.220 156.470 121.290 ;
        RECT 134.980 119.710 135.150 121.120 ;
        RECT 135.490 120.250 135.660 120.580 ;
        RECT 135.875 120.550 136.915 120.720 ;
        RECT 135.875 120.110 136.915 120.280 ;
        RECT 137.130 120.250 137.300 120.580 ;
        RECT 137.640 119.710 137.930 121.120 ;
        RECT 134.980 119.590 137.930 119.710 ;
        RECT 153.600 121.120 156.470 121.220 ;
        RECT 153.600 119.710 153.900 121.120 ;
        RECT 154.240 120.250 154.410 120.580 ;
        RECT 154.580 120.550 155.620 120.720 ;
        RECT 154.580 120.110 155.620 120.280 ;
        RECT 155.790 120.250 155.960 120.580 ;
        RECT 156.300 119.710 156.470 121.120 ;
        RECT 134.980 119.540 137.810 119.590 ;
        RECT 153.600 119.570 156.470 119.710 ;
        RECT 153.730 119.540 156.470 119.570 ;
        RECT 157.030 121.250 159.860 121.300 ;
        RECT 157.030 121.130 159.980 121.250 ;
        RECT 157.030 119.720 157.200 121.130 ;
        RECT 157.540 120.260 157.710 120.590 ;
        RECT 157.925 120.560 158.965 120.730 ;
        RECT 157.925 120.120 158.965 120.290 ;
        RECT 159.180 120.260 159.350 120.590 ;
        RECT 159.690 119.720 159.980 121.130 ;
        RECT 157.030 119.600 159.980 119.720 ;
        RECT 157.030 119.550 159.860 119.600 ;
        RECT 131.680 119.110 134.420 119.180 ;
        RECT 131.550 119.010 134.420 119.110 ;
        RECT 131.550 117.600 131.850 119.010 ;
        RECT 132.190 118.140 132.360 118.470 ;
        RECT 132.530 118.440 133.570 118.610 ;
        RECT 132.530 118.000 133.570 118.170 ;
        RECT 133.740 118.140 133.910 118.470 ;
        RECT 134.250 117.600 134.420 119.010 ;
        RECT 131.550 117.460 134.420 117.600 ;
        RECT 131.680 117.430 134.420 117.460 ;
        RECT 134.980 119.140 137.810 119.190 ;
        RECT 134.980 119.020 137.930 119.140 ;
        RECT 153.730 119.120 156.470 119.190 ;
        RECT 134.980 117.610 135.150 119.020 ;
        RECT 135.490 118.150 135.660 118.480 ;
        RECT 135.875 118.450 136.915 118.620 ;
        RECT 135.875 118.010 136.915 118.180 ;
        RECT 137.130 118.150 137.300 118.480 ;
        RECT 137.640 117.610 137.930 119.020 ;
        RECT 134.980 117.490 137.930 117.610 ;
        RECT 153.600 119.020 156.470 119.120 ;
        RECT 153.600 117.610 153.900 119.020 ;
        RECT 154.240 118.150 154.410 118.480 ;
        RECT 154.580 118.450 155.620 118.620 ;
        RECT 154.580 118.010 155.620 118.180 ;
        RECT 155.790 118.150 155.960 118.480 ;
        RECT 156.300 117.610 156.470 119.020 ;
        RECT 134.980 117.440 137.810 117.490 ;
        RECT 153.600 117.470 156.470 117.610 ;
        RECT 153.730 117.440 156.470 117.470 ;
        RECT 157.030 119.150 159.860 119.200 ;
        RECT 157.030 119.030 159.980 119.150 ;
        RECT 157.030 117.620 157.200 119.030 ;
        RECT 157.540 118.160 157.710 118.490 ;
        RECT 157.925 118.460 158.965 118.630 ;
        RECT 157.925 118.020 158.965 118.190 ;
        RECT 159.180 118.160 159.350 118.490 ;
        RECT 159.690 117.620 159.980 119.030 ;
        RECT 157.030 117.500 159.980 117.620 ;
        RECT 157.030 117.450 159.860 117.500 ;
        RECT 131.680 117.010 134.420 117.080 ;
        RECT 131.550 116.910 134.420 117.010 ;
        RECT 131.550 115.500 131.850 116.910 ;
        RECT 132.190 116.040 132.360 116.370 ;
        RECT 132.530 116.340 133.570 116.510 ;
        RECT 132.530 115.900 133.570 116.070 ;
        RECT 133.740 116.040 133.910 116.370 ;
        RECT 134.250 115.500 134.420 116.910 ;
        RECT 131.550 115.360 134.420 115.500 ;
        RECT 131.680 115.330 134.420 115.360 ;
        RECT 134.980 117.040 137.810 117.090 ;
        RECT 134.980 116.920 137.930 117.040 ;
        RECT 153.730 117.020 156.470 117.090 ;
        RECT 134.980 115.510 135.150 116.920 ;
        RECT 135.490 116.050 135.660 116.380 ;
        RECT 135.875 116.350 136.915 116.520 ;
        RECT 135.875 115.910 136.915 116.080 ;
        RECT 137.130 116.050 137.300 116.380 ;
        RECT 137.640 115.510 137.930 116.920 ;
        RECT 134.980 115.390 137.930 115.510 ;
        RECT 153.600 116.920 156.470 117.020 ;
        RECT 153.600 115.510 153.900 116.920 ;
        RECT 154.240 116.050 154.410 116.380 ;
        RECT 154.580 116.350 155.620 116.520 ;
        RECT 154.580 115.910 155.620 116.080 ;
        RECT 155.790 116.050 155.960 116.380 ;
        RECT 156.300 115.510 156.470 116.920 ;
        RECT 134.980 115.340 137.810 115.390 ;
        RECT 153.600 115.370 156.470 115.510 ;
        RECT 153.730 115.340 156.470 115.370 ;
        RECT 157.030 117.050 159.860 117.100 ;
        RECT 157.030 116.930 159.980 117.050 ;
        RECT 157.030 115.520 157.200 116.930 ;
        RECT 157.540 116.060 157.710 116.390 ;
        RECT 157.925 116.360 158.965 116.530 ;
        RECT 157.925 115.920 158.965 116.090 ;
        RECT 159.180 116.060 159.350 116.390 ;
        RECT 159.690 115.520 159.980 116.930 ;
        RECT 157.030 115.400 159.980 115.520 ;
        RECT 157.030 115.350 159.860 115.400 ;
        RECT 131.680 114.910 134.420 114.980 ;
        RECT 131.550 114.810 134.420 114.910 ;
        RECT 131.550 113.400 131.850 114.810 ;
        RECT 132.190 113.940 132.360 114.270 ;
        RECT 132.530 114.240 133.570 114.410 ;
        RECT 132.530 113.800 133.570 113.970 ;
        RECT 133.740 113.940 133.910 114.270 ;
        RECT 134.250 113.400 134.420 114.810 ;
        RECT 131.550 113.260 134.420 113.400 ;
        RECT 131.680 113.230 134.420 113.260 ;
        RECT 134.980 114.940 137.810 114.990 ;
        RECT 134.980 114.820 137.930 114.940 ;
        RECT 153.730 114.920 156.470 114.990 ;
        RECT 134.980 113.410 135.150 114.820 ;
        RECT 135.490 113.950 135.660 114.280 ;
        RECT 135.875 114.250 136.915 114.420 ;
        RECT 135.875 113.810 136.915 113.980 ;
        RECT 137.130 113.950 137.300 114.280 ;
        RECT 137.640 113.410 137.930 114.820 ;
        RECT 134.980 113.290 137.930 113.410 ;
        RECT 153.600 114.820 156.470 114.920 ;
        RECT 153.600 113.410 153.900 114.820 ;
        RECT 154.240 113.950 154.410 114.280 ;
        RECT 154.580 114.250 155.620 114.420 ;
        RECT 154.580 113.810 155.620 113.980 ;
        RECT 155.790 113.950 155.960 114.280 ;
        RECT 156.300 113.410 156.470 114.820 ;
        RECT 134.980 113.240 137.810 113.290 ;
        RECT 153.600 113.270 156.470 113.410 ;
        RECT 153.730 113.240 156.470 113.270 ;
        RECT 157.030 114.950 159.860 115.000 ;
        RECT 157.030 114.830 159.980 114.950 ;
        RECT 157.030 113.420 157.200 114.830 ;
        RECT 157.540 113.960 157.710 114.290 ;
        RECT 157.925 114.260 158.965 114.430 ;
        RECT 157.925 113.820 158.965 113.990 ;
        RECT 159.180 113.960 159.350 114.290 ;
        RECT 159.690 113.420 159.980 114.830 ;
        RECT 157.030 113.300 159.980 113.420 ;
        RECT 157.030 113.250 159.860 113.300 ;
        RECT 131.680 112.810 134.420 112.880 ;
        RECT 131.550 112.710 134.420 112.810 ;
        RECT 131.550 111.300 131.850 112.710 ;
        RECT 132.190 111.840 132.360 112.170 ;
        RECT 132.530 112.140 133.570 112.310 ;
        RECT 132.530 111.700 133.570 111.870 ;
        RECT 133.740 111.840 133.910 112.170 ;
        RECT 134.250 111.300 134.420 112.710 ;
        RECT 131.550 111.160 134.420 111.300 ;
        RECT 131.680 111.130 134.420 111.160 ;
        RECT 134.980 112.840 137.810 112.890 ;
        RECT 134.980 112.720 137.930 112.840 ;
        RECT 153.730 112.820 156.470 112.890 ;
        RECT 134.980 111.310 135.150 112.720 ;
        RECT 135.490 111.850 135.660 112.180 ;
        RECT 135.875 112.150 136.915 112.320 ;
        RECT 135.875 111.710 136.915 111.880 ;
        RECT 137.130 111.850 137.300 112.180 ;
        RECT 137.640 111.310 137.930 112.720 ;
        RECT 134.980 111.190 137.930 111.310 ;
        RECT 153.600 112.720 156.470 112.820 ;
        RECT 153.600 111.310 153.900 112.720 ;
        RECT 154.240 111.850 154.410 112.180 ;
        RECT 154.580 112.150 155.620 112.320 ;
        RECT 154.580 111.710 155.620 111.880 ;
        RECT 155.790 111.850 155.960 112.180 ;
        RECT 156.300 111.310 156.470 112.720 ;
        RECT 134.980 111.140 137.810 111.190 ;
        RECT 153.600 111.170 156.470 111.310 ;
        RECT 153.730 111.140 156.470 111.170 ;
        RECT 157.030 112.850 159.860 112.900 ;
        RECT 157.030 112.730 159.980 112.850 ;
        RECT 157.030 111.320 157.200 112.730 ;
        RECT 157.540 111.860 157.710 112.190 ;
        RECT 157.925 112.160 158.965 112.330 ;
        RECT 157.925 111.720 158.965 111.890 ;
        RECT 159.180 111.860 159.350 112.190 ;
        RECT 159.690 111.320 159.980 112.730 ;
        RECT 157.030 111.200 159.980 111.320 ;
        RECT 157.030 111.150 159.860 111.200 ;
        RECT 131.680 110.710 134.420 110.780 ;
        RECT 131.550 110.610 134.420 110.710 ;
        RECT 131.550 109.200 131.850 110.610 ;
        RECT 132.190 109.740 132.360 110.070 ;
        RECT 132.530 110.040 133.570 110.210 ;
        RECT 132.530 109.600 133.570 109.770 ;
        RECT 133.740 109.740 133.910 110.070 ;
        RECT 134.250 109.200 134.420 110.610 ;
        RECT 131.550 109.060 134.420 109.200 ;
        RECT 131.680 109.030 134.420 109.060 ;
        RECT 134.980 110.740 137.810 110.790 ;
        RECT 134.980 110.620 137.930 110.740 ;
        RECT 153.730 110.720 156.470 110.790 ;
        RECT 134.980 109.210 135.150 110.620 ;
        RECT 135.490 109.750 135.660 110.080 ;
        RECT 135.875 110.050 136.915 110.220 ;
        RECT 135.875 109.610 136.915 109.780 ;
        RECT 137.130 109.750 137.300 110.080 ;
        RECT 137.640 109.210 137.930 110.620 ;
        RECT 134.980 109.090 137.930 109.210 ;
        RECT 153.600 110.620 156.470 110.720 ;
        RECT 153.600 109.210 153.900 110.620 ;
        RECT 154.240 109.750 154.410 110.080 ;
        RECT 154.580 110.050 155.620 110.220 ;
        RECT 154.580 109.610 155.620 109.780 ;
        RECT 155.790 109.750 155.960 110.080 ;
        RECT 156.300 109.210 156.470 110.620 ;
        RECT 134.980 109.040 137.810 109.090 ;
        RECT 153.600 109.070 156.470 109.210 ;
        RECT 153.730 109.040 156.470 109.070 ;
        RECT 157.030 110.750 159.860 110.800 ;
        RECT 157.030 110.630 159.980 110.750 ;
        RECT 157.030 109.220 157.200 110.630 ;
        RECT 157.540 109.760 157.710 110.090 ;
        RECT 157.925 110.060 158.965 110.230 ;
        RECT 157.925 109.620 158.965 109.790 ;
        RECT 159.180 109.760 159.350 110.090 ;
        RECT 159.690 109.220 159.980 110.630 ;
        RECT 157.030 109.100 159.980 109.220 ;
        RECT 157.030 109.050 159.860 109.100 ;
        RECT 131.680 108.610 134.420 108.680 ;
        RECT 131.550 108.510 134.420 108.610 ;
        RECT 131.550 107.100 131.850 108.510 ;
        RECT 132.190 107.640 132.360 107.970 ;
        RECT 132.530 107.940 133.570 108.110 ;
        RECT 132.530 107.500 133.570 107.670 ;
        RECT 133.740 107.640 133.910 107.970 ;
        RECT 134.250 107.100 134.420 108.510 ;
        RECT 131.550 106.960 134.420 107.100 ;
        RECT 131.680 106.930 134.420 106.960 ;
        RECT 134.980 108.640 137.810 108.690 ;
        RECT 134.980 108.520 137.930 108.640 ;
        RECT 153.730 108.620 156.470 108.690 ;
        RECT 134.980 107.110 135.150 108.520 ;
        RECT 135.490 107.650 135.660 107.980 ;
        RECT 135.875 107.950 136.915 108.120 ;
        RECT 135.875 107.510 136.915 107.680 ;
        RECT 137.130 107.650 137.300 107.980 ;
        RECT 137.640 107.110 137.930 108.520 ;
        RECT 134.980 106.990 137.930 107.110 ;
        RECT 153.600 108.520 156.470 108.620 ;
        RECT 153.600 107.110 153.900 108.520 ;
        RECT 154.240 107.650 154.410 107.980 ;
        RECT 154.580 107.950 155.620 108.120 ;
        RECT 154.580 107.510 155.620 107.680 ;
        RECT 155.790 107.650 155.960 107.980 ;
        RECT 156.300 107.110 156.470 108.520 ;
        RECT 134.980 106.940 137.810 106.990 ;
        RECT 153.600 106.970 156.470 107.110 ;
        RECT 153.730 106.940 156.470 106.970 ;
        RECT 157.030 108.650 159.860 108.700 ;
        RECT 157.030 108.530 159.980 108.650 ;
        RECT 157.030 107.120 157.200 108.530 ;
        RECT 157.540 107.660 157.710 107.990 ;
        RECT 157.925 107.960 158.965 108.130 ;
        RECT 157.925 107.520 158.965 107.690 ;
        RECT 159.180 107.660 159.350 107.990 ;
        RECT 159.690 107.120 159.980 108.530 ;
        RECT 157.030 107.000 159.980 107.120 ;
        RECT 157.030 106.950 159.860 107.000 ;
        RECT 131.680 106.510 134.420 106.580 ;
        RECT 131.550 106.410 134.420 106.510 ;
        RECT 131.550 105.000 131.850 106.410 ;
        RECT 132.190 105.540 132.360 105.870 ;
        RECT 132.530 105.840 133.570 106.010 ;
        RECT 132.530 105.400 133.570 105.570 ;
        RECT 133.740 105.540 133.910 105.870 ;
        RECT 134.250 105.000 134.420 106.410 ;
        RECT 131.550 104.860 134.420 105.000 ;
        RECT 131.680 104.830 134.420 104.860 ;
        RECT 134.980 106.540 137.810 106.590 ;
        RECT 134.980 106.420 137.930 106.540 ;
        RECT 153.730 106.520 156.470 106.590 ;
        RECT 134.980 105.010 135.150 106.420 ;
        RECT 135.490 105.550 135.660 105.880 ;
        RECT 135.875 105.850 136.915 106.020 ;
        RECT 135.875 105.410 136.915 105.580 ;
        RECT 137.130 105.550 137.300 105.880 ;
        RECT 137.640 105.010 137.930 106.420 ;
        RECT 134.980 104.890 137.930 105.010 ;
        RECT 153.600 106.420 156.470 106.520 ;
        RECT 153.600 105.010 153.900 106.420 ;
        RECT 154.240 105.550 154.410 105.880 ;
        RECT 154.580 105.850 155.620 106.020 ;
        RECT 154.580 105.410 155.620 105.580 ;
        RECT 155.790 105.550 155.960 105.880 ;
        RECT 156.300 105.010 156.470 106.420 ;
        RECT 134.980 104.840 137.810 104.890 ;
        RECT 153.600 104.870 156.470 105.010 ;
        RECT 153.730 104.840 156.470 104.870 ;
        RECT 157.030 106.550 159.860 106.600 ;
        RECT 157.030 106.430 159.980 106.550 ;
        RECT 157.030 105.020 157.200 106.430 ;
        RECT 157.540 105.560 157.710 105.890 ;
        RECT 157.925 105.860 158.965 106.030 ;
        RECT 157.925 105.420 158.965 105.590 ;
        RECT 159.180 105.560 159.350 105.890 ;
        RECT 159.690 105.020 159.980 106.430 ;
        RECT 157.030 104.900 159.980 105.020 ;
        RECT 157.030 104.850 159.860 104.900 ;
        RECT 131.680 104.410 134.420 104.480 ;
        RECT 131.550 104.310 134.420 104.410 ;
        RECT 131.550 102.900 131.850 104.310 ;
        RECT 132.190 103.440 132.360 103.770 ;
        RECT 132.530 103.740 133.570 103.910 ;
        RECT 132.530 103.300 133.570 103.470 ;
        RECT 133.740 103.440 133.910 103.770 ;
        RECT 134.250 102.900 134.420 104.310 ;
        RECT 131.550 102.760 134.420 102.900 ;
        RECT 131.680 102.730 134.420 102.760 ;
        RECT 134.980 104.440 137.810 104.490 ;
        RECT 134.980 104.320 137.930 104.440 ;
        RECT 153.730 104.420 156.470 104.490 ;
        RECT 134.980 102.910 135.150 104.320 ;
        RECT 135.490 103.450 135.660 103.780 ;
        RECT 135.875 103.750 136.915 103.920 ;
        RECT 135.875 103.310 136.915 103.480 ;
        RECT 137.130 103.450 137.300 103.780 ;
        RECT 137.640 102.910 137.930 104.320 ;
        RECT 134.980 102.790 137.930 102.910 ;
        RECT 153.600 104.320 156.470 104.420 ;
        RECT 153.600 102.910 153.900 104.320 ;
        RECT 154.240 103.450 154.410 103.780 ;
        RECT 154.580 103.750 155.620 103.920 ;
        RECT 154.580 103.310 155.620 103.480 ;
        RECT 155.790 103.450 155.960 103.780 ;
        RECT 156.300 102.910 156.470 104.320 ;
        RECT 134.980 102.740 137.810 102.790 ;
        RECT 153.600 102.770 156.470 102.910 ;
        RECT 153.730 102.740 156.470 102.770 ;
        RECT 157.030 104.450 159.860 104.500 ;
        RECT 157.030 104.330 159.980 104.450 ;
        RECT 157.030 102.920 157.200 104.330 ;
        RECT 157.540 103.460 157.710 103.790 ;
        RECT 157.925 103.760 158.965 103.930 ;
        RECT 157.925 103.320 158.965 103.490 ;
        RECT 159.180 103.460 159.350 103.790 ;
        RECT 159.690 102.920 159.980 104.330 ;
        RECT 157.030 102.800 159.980 102.920 ;
        RECT 157.030 102.750 159.860 102.800 ;
        RECT 131.680 102.310 134.420 102.380 ;
        RECT 131.550 102.210 134.420 102.310 ;
        RECT 131.550 100.800 131.850 102.210 ;
        RECT 132.190 101.340 132.360 101.670 ;
        RECT 132.530 101.640 133.570 101.810 ;
        RECT 132.530 101.200 133.570 101.370 ;
        RECT 133.740 101.340 133.910 101.670 ;
        RECT 134.250 100.800 134.420 102.210 ;
        RECT 131.550 100.660 134.420 100.800 ;
        RECT 131.680 100.630 134.420 100.660 ;
        RECT 134.980 102.340 137.810 102.390 ;
        RECT 134.980 102.220 137.930 102.340 ;
        RECT 153.730 102.320 156.470 102.390 ;
        RECT 134.980 100.810 135.150 102.220 ;
        RECT 135.490 101.350 135.660 101.680 ;
        RECT 135.875 101.650 136.915 101.820 ;
        RECT 135.875 101.210 136.915 101.380 ;
        RECT 137.130 101.350 137.300 101.680 ;
        RECT 137.640 100.810 137.930 102.220 ;
        RECT 134.980 100.690 137.930 100.810 ;
        RECT 153.600 102.220 156.470 102.320 ;
        RECT 153.600 100.810 153.900 102.220 ;
        RECT 154.240 101.350 154.410 101.680 ;
        RECT 154.580 101.650 155.620 101.820 ;
        RECT 154.580 101.210 155.620 101.380 ;
        RECT 155.790 101.350 155.960 101.680 ;
        RECT 156.300 100.810 156.470 102.220 ;
        RECT 134.980 100.640 137.810 100.690 ;
        RECT 153.600 100.670 156.470 100.810 ;
        RECT 153.730 100.640 156.470 100.670 ;
        RECT 157.030 102.350 159.860 102.400 ;
        RECT 157.030 102.230 159.980 102.350 ;
        RECT 157.030 100.820 157.200 102.230 ;
        RECT 157.540 101.360 157.710 101.690 ;
        RECT 157.925 101.660 158.965 101.830 ;
        RECT 157.925 101.220 158.965 101.390 ;
        RECT 159.180 101.360 159.350 101.690 ;
        RECT 159.690 100.820 159.980 102.230 ;
        RECT 157.030 100.700 159.980 100.820 ;
        RECT 157.030 100.650 159.860 100.700 ;
        RECT 131.680 100.210 134.420 100.280 ;
        RECT 131.550 100.110 134.420 100.210 ;
        RECT 131.550 98.700 131.850 100.110 ;
        RECT 132.190 99.240 132.360 99.570 ;
        RECT 132.530 99.540 133.570 99.710 ;
        RECT 132.530 99.100 133.570 99.270 ;
        RECT 133.740 99.240 133.910 99.570 ;
        RECT 134.250 98.700 134.420 100.110 ;
        RECT 131.550 98.560 134.420 98.700 ;
        RECT 131.680 98.530 134.420 98.560 ;
        RECT 134.980 100.240 137.810 100.290 ;
        RECT 134.980 100.120 137.930 100.240 ;
        RECT 153.730 100.220 156.470 100.290 ;
        RECT 134.980 98.710 135.150 100.120 ;
        RECT 135.490 99.250 135.660 99.580 ;
        RECT 135.875 99.550 136.915 99.720 ;
        RECT 135.875 99.110 136.915 99.280 ;
        RECT 137.130 99.250 137.300 99.580 ;
        RECT 137.640 98.710 137.930 100.120 ;
        RECT 134.980 98.590 137.930 98.710 ;
        RECT 153.600 100.120 156.470 100.220 ;
        RECT 153.600 98.710 153.900 100.120 ;
        RECT 154.240 99.250 154.410 99.580 ;
        RECT 154.580 99.550 155.620 99.720 ;
        RECT 154.580 99.110 155.620 99.280 ;
        RECT 155.790 99.250 155.960 99.580 ;
        RECT 156.300 98.710 156.470 100.120 ;
        RECT 134.980 98.540 137.810 98.590 ;
        RECT 153.600 98.570 156.470 98.710 ;
        RECT 153.730 98.540 156.470 98.570 ;
        RECT 157.030 100.250 159.860 100.300 ;
        RECT 157.030 100.130 159.980 100.250 ;
        RECT 157.030 98.720 157.200 100.130 ;
        RECT 157.540 99.260 157.710 99.590 ;
        RECT 157.925 99.560 158.965 99.730 ;
        RECT 157.925 99.120 158.965 99.290 ;
        RECT 159.180 99.260 159.350 99.590 ;
        RECT 159.690 98.720 159.980 100.130 ;
        RECT 157.030 98.600 159.980 98.720 ;
        RECT 157.030 98.550 159.860 98.600 ;
        RECT 131.680 98.110 134.420 98.180 ;
        RECT 131.550 98.010 134.420 98.110 ;
        RECT 131.550 96.600 131.850 98.010 ;
        RECT 132.190 97.140 132.360 97.470 ;
        RECT 132.530 97.440 133.570 97.610 ;
        RECT 132.530 97.000 133.570 97.170 ;
        RECT 133.740 97.140 133.910 97.470 ;
        RECT 134.250 96.600 134.420 98.010 ;
        RECT 131.550 96.460 134.420 96.600 ;
        RECT 131.680 96.430 134.420 96.460 ;
        RECT 134.980 98.140 137.810 98.190 ;
        RECT 134.980 98.020 137.930 98.140 ;
        RECT 153.730 98.120 156.470 98.190 ;
        RECT 134.980 96.610 135.150 98.020 ;
        RECT 135.490 97.150 135.660 97.480 ;
        RECT 135.875 97.450 136.915 97.620 ;
        RECT 135.875 97.010 136.915 97.180 ;
        RECT 137.130 97.150 137.300 97.480 ;
        RECT 137.640 96.610 137.930 98.020 ;
        RECT 134.980 96.490 137.930 96.610 ;
        RECT 153.600 98.020 156.470 98.120 ;
        RECT 153.600 96.610 153.900 98.020 ;
        RECT 154.240 97.150 154.410 97.480 ;
        RECT 154.580 97.450 155.620 97.620 ;
        RECT 154.580 97.010 155.620 97.180 ;
        RECT 155.790 97.150 155.960 97.480 ;
        RECT 156.300 96.610 156.470 98.020 ;
        RECT 134.980 96.440 137.810 96.490 ;
        RECT 153.600 96.470 156.470 96.610 ;
        RECT 153.730 96.440 156.470 96.470 ;
        RECT 157.030 98.150 159.860 98.200 ;
        RECT 157.030 98.030 159.980 98.150 ;
        RECT 157.030 96.620 157.200 98.030 ;
        RECT 157.540 97.160 157.710 97.490 ;
        RECT 157.925 97.460 158.965 97.630 ;
        RECT 157.925 97.020 158.965 97.190 ;
        RECT 159.180 97.160 159.350 97.490 ;
        RECT 159.690 96.620 159.980 98.030 ;
        RECT 157.030 96.500 159.980 96.620 ;
        RECT 157.030 96.450 159.860 96.500 ;
        RECT 131.680 96.010 134.420 96.080 ;
        RECT 131.550 95.910 134.420 96.010 ;
        RECT 131.550 94.500 131.850 95.910 ;
        RECT 132.190 95.040 132.360 95.370 ;
        RECT 132.530 95.340 133.570 95.510 ;
        RECT 132.530 94.900 133.570 95.070 ;
        RECT 133.740 95.040 133.910 95.370 ;
        RECT 134.250 94.500 134.420 95.910 ;
        RECT 131.550 94.360 134.420 94.500 ;
        RECT 131.680 94.330 134.420 94.360 ;
        RECT 134.980 96.040 137.810 96.090 ;
        RECT 134.980 95.920 137.930 96.040 ;
        RECT 153.730 96.020 156.470 96.090 ;
        RECT 134.980 94.510 135.150 95.920 ;
        RECT 135.490 95.050 135.660 95.380 ;
        RECT 135.875 95.350 136.915 95.520 ;
        RECT 135.875 94.910 136.915 95.080 ;
        RECT 137.130 95.050 137.300 95.380 ;
        RECT 137.640 94.510 137.930 95.920 ;
        RECT 134.980 94.390 137.930 94.510 ;
        RECT 153.600 95.920 156.470 96.020 ;
        RECT 153.600 94.510 153.900 95.920 ;
        RECT 154.240 95.050 154.410 95.380 ;
        RECT 154.580 95.350 155.620 95.520 ;
        RECT 154.580 94.910 155.620 95.080 ;
        RECT 155.790 95.050 155.960 95.380 ;
        RECT 156.300 94.510 156.470 95.920 ;
        RECT 134.980 94.340 137.810 94.390 ;
        RECT 153.600 94.370 156.470 94.510 ;
        RECT 153.730 94.340 156.470 94.370 ;
        RECT 157.030 96.050 159.860 96.100 ;
        RECT 157.030 95.930 159.980 96.050 ;
        RECT 157.030 94.520 157.200 95.930 ;
        RECT 157.540 95.060 157.710 95.390 ;
        RECT 157.925 95.360 158.965 95.530 ;
        RECT 157.925 94.920 158.965 95.090 ;
        RECT 159.180 95.060 159.350 95.390 ;
        RECT 159.690 94.520 159.980 95.930 ;
        RECT 157.030 94.400 159.980 94.520 ;
        RECT 157.030 94.350 159.860 94.400 ;
        RECT 131.680 93.910 134.420 93.980 ;
        RECT 131.550 93.810 134.420 93.910 ;
        RECT 131.550 92.400 131.850 93.810 ;
        RECT 132.190 92.940 132.360 93.270 ;
        RECT 132.530 93.240 133.570 93.410 ;
        RECT 132.530 92.800 133.570 92.970 ;
        RECT 133.740 92.940 133.910 93.270 ;
        RECT 134.250 92.400 134.420 93.810 ;
        RECT 131.550 92.260 134.420 92.400 ;
        RECT 131.680 92.230 134.420 92.260 ;
        RECT 134.980 93.940 137.810 93.990 ;
        RECT 134.980 93.820 137.930 93.940 ;
        RECT 153.730 93.920 156.470 93.990 ;
        RECT 134.980 92.410 135.150 93.820 ;
        RECT 135.490 92.950 135.660 93.280 ;
        RECT 135.875 93.250 136.915 93.420 ;
        RECT 135.875 92.810 136.915 92.980 ;
        RECT 137.130 92.950 137.300 93.280 ;
        RECT 137.640 92.410 137.930 93.820 ;
        RECT 134.980 92.290 137.930 92.410 ;
        RECT 153.600 93.820 156.470 93.920 ;
        RECT 153.600 92.410 153.900 93.820 ;
        RECT 154.240 92.950 154.410 93.280 ;
        RECT 154.580 93.250 155.620 93.420 ;
        RECT 154.580 92.810 155.620 92.980 ;
        RECT 155.790 92.950 155.960 93.280 ;
        RECT 156.300 92.410 156.470 93.820 ;
        RECT 134.980 92.240 137.810 92.290 ;
        RECT 153.600 92.270 156.470 92.410 ;
        RECT 153.730 92.240 156.470 92.270 ;
        RECT 157.030 93.950 159.860 94.000 ;
        RECT 157.030 93.830 159.980 93.950 ;
        RECT 157.030 92.420 157.200 93.830 ;
        RECT 157.540 92.960 157.710 93.290 ;
        RECT 157.925 93.260 158.965 93.430 ;
        RECT 157.925 92.820 158.965 92.990 ;
        RECT 159.180 92.960 159.350 93.290 ;
        RECT 159.690 92.420 159.980 93.830 ;
        RECT 157.030 92.300 159.980 92.420 ;
        RECT 157.030 92.250 159.860 92.300 ;
        RECT 131.680 91.810 134.420 91.880 ;
        RECT 131.550 91.710 134.420 91.810 ;
        RECT 131.550 90.300 131.850 91.710 ;
        RECT 132.190 90.840 132.360 91.170 ;
        RECT 132.530 91.140 133.570 91.310 ;
        RECT 132.530 90.700 133.570 90.870 ;
        RECT 133.740 90.840 133.910 91.170 ;
        RECT 134.250 90.300 134.420 91.710 ;
        RECT 131.550 90.160 134.420 90.300 ;
        RECT 131.680 90.130 134.420 90.160 ;
        RECT 134.980 91.840 137.810 91.890 ;
        RECT 134.980 91.720 137.930 91.840 ;
        RECT 153.730 91.820 156.470 91.890 ;
        RECT 134.980 90.310 135.150 91.720 ;
        RECT 135.490 90.850 135.660 91.180 ;
        RECT 135.875 91.150 136.915 91.320 ;
        RECT 135.875 90.710 136.915 90.880 ;
        RECT 137.130 90.850 137.300 91.180 ;
        RECT 137.640 90.310 137.930 91.720 ;
        RECT 134.980 90.190 137.930 90.310 ;
        RECT 153.600 91.720 156.470 91.820 ;
        RECT 153.600 90.310 153.900 91.720 ;
        RECT 154.240 90.850 154.410 91.180 ;
        RECT 154.580 91.150 155.620 91.320 ;
        RECT 154.580 90.710 155.620 90.880 ;
        RECT 155.790 90.850 155.960 91.180 ;
        RECT 156.300 90.310 156.470 91.720 ;
        RECT 134.980 90.140 137.810 90.190 ;
        RECT 153.600 90.170 156.470 90.310 ;
        RECT 153.730 90.140 156.470 90.170 ;
        RECT 157.030 91.850 159.860 91.900 ;
        RECT 157.030 91.730 159.980 91.850 ;
        RECT 157.030 90.320 157.200 91.730 ;
        RECT 157.540 90.860 157.710 91.190 ;
        RECT 157.925 91.160 158.965 91.330 ;
        RECT 157.925 90.720 158.965 90.890 ;
        RECT 159.180 90.860 159.350 91.190 ;
        RECT 159.690 90.320 159.980 91.730 ;
        RECT 157.030 90.200 159.980 90.320 ;
        RECT 157.030 90.150 159.860 90.200 ;
        RECT 131.680 89.710 134.420 89.780 ;
        RECT 131.550 89.610 134.420 89.710 ;
        RECT 131.550 88.200 131.850 89.610 ;
        RECT 132.190 88.740 132.360 89.070 ;
        RECT 132.530 89.040 133.570 89.210 ;
        RECT 132.530 88.600 133.570 88.770 ;
        RECT 133.740 88.740 133.910 89.070 ;
        RECT 134.250 88.200 134.420 89.610 ;
        RECT 131.550 88.060 134.420 88.200 ;
        RECT 131.680 88.030 134.420 88.060 ;
        RECT 134.980 89.740 137.810 89.790 ;
        RECT 134.980 89.620 137.930 89.740 ;
        RECT 153.730 89.720 156.470 89.790 ;
        RECT 134.980 88.210 135.150 89.620 ;
        RECT 135.490 88.750 135.660 89.080 ;
        RECT 135.875 89.050 136.915 89.220 ;
        RECT 135.875 88.610 136.915 88.780 ;
        RECT 137.130 88.750 137.300 89.080 ;
        RECT 137.640 88.210 137.930 89.620 ;
        RECT 134.980 88.090 137.930 88.210 ;
        RECT 153.600 89.620 156.470 89.720 ;
        RECT 153.600 88.210 153.900 89.620 ;
        RECT 154.240 88.750 154.410 89.080 ;
        RECT 154.580 89.050 155.620 89.220 ;
        RECT 154.580 88.610 155.620 88.780 ;
        RECT 155.790 88.750 155.960 89.080 ;
        RECT 156.300 88.210 156.470 89.620 ;
        RECT 134.980 88.040 137.810 88.090 ;
        RECT 153.600 88.070 156.470 88.210 ;
        RECT 153.730 88.040 156.470 88.070 ;
        RECT 157.030 89.750 159.860 89.800 ;
        RECT 157.030 89.630 159.980 89.750 ;
        RECT 157.030 88.220 157.200 89.630 ;
        RECT 157.540 88.760 157.710 89.090 ;
        RECT 157.925 89.060 158.965 89.230 ;
        RECT 157.925 88.620 158.965 88.790 ;
        RECT 159.180 88.760 159.350 89.090 ;
        RECT 159.690 88.220 159.980 89.630 ;
        RECT 157.030 88.100 159.980 88.220 ;
        RECT 157.030 88.050 159.860 88.100 ;
        RECT 131.680 87.610 134.420 87.680 ;
        RECT 131.550 87.510 134.420 87.610 ;
        RECT 131.550 86.100 131.850 87.510 ;
        RECT 132.190 86.640 132.360 86.970 ;
        RECT 132.530 86.940 133.570 87.110 ;
        RECT 132.530 86.500 133.570 86.670 ;
        RECT 133.740 86.640 133.910 86.970 ;
        RECT 134.250 86.100 134.420 87.510 ;
        RECT 131.550 85.960 134.420 86.100 ;
        RECT 131.680 85.930 134.420 85.960 ;
        RECT 134.980 87.640 137.810 87.690 ;
        RECT 134.980 87.520 137.930 87.640 ;
        RECT 153.730 87.620 156.470 87.690 ;
        RECT 134.980 86.110 135.150 87.520 ;
        RECT 135.490 86.650 135.660 86.980 ;
        RECT 135.875 86.950 136.915 87.120 ;
        RECT 135.875 86.510 136.915 86.680 ;
        RECT 137.130 86.650 137.300 86.980 ;
        RECT 137.640 86.110 137.930 87.520 ;
        RECT 134.980 85.990 137.930 86.110 ;
        RECT 153.600 87.520 156.470 87.620 ;
        RECT 153.600 86.110 153.900 87.520 ;
        RECT 154.240 86.650 154.410 86.980 ;
        RECT 154.580 86.950 155.620 87.120 ;
        RECT 154.580 86.510 155.620 86.680 ;
        RECT 155.790 86.650 155.960 86.980 ;
        RECT 156.300 86.110 156.470 87.520 ;
        RECT 134.980 85.940 137.810 85.990 ;
        RECT 153.600 85.970 156.470 86.110 ;
        RECT 153.730 85.940 156.470 85.970 ;
        RECT 157.030 87.650 159.860 87.700 ;
        RECT 157.030 87.530 159.980 87.650 ;
        RECT 157.030 86.120 157.200 87.530 ;
        RECT 157.540 86.660 157.710 86.990 ;
        RECT 157.925 86.960 158.965 87.130 ;
        RECT 157.925 86.520 158.965 86.690 ;
        RECT 159.180 86.660 159.350 86.990 ;
        RECT 159.690 86.120 159.980 87.530 ;
        RECT 157.030 86.000 159.980 86.120 ;
        RECT 157.030 85.950 159.860 86.000 ;
        RECT 131.680 85.510 134.420 85.580 ;
        RECT 131.550 85.410 134.420 85.510 ;
        RECT 131.550 84.000 131.850 85.410 ;
        RECT 132.190 84.540 132.360 84.870 ;
        RECT 132.530 84.840 133.570 85.010 ;
        RECT 132.530 84.400 133.570 84.570 ;
        RECT 133.740 84.540 133.910 84.870 ;
        RECT 134.250 84.000 134.420 85.410 ;
        RECT 131.550 83.860 134.420 84.000 ;
        RECT 131.680 83.830 134.420 83.860 ;
        RECT 134.980 85.540 137.810 85.590 ;
        RECT 134.980 85.420 137.930 85.540 ;
        RECT 153.730 85.520 156.470 85.590 ;
        RECT 134.980 84.010 135.150 85.420 ;
        RECT 135.490 84.550 135.660 84.880 ;
        RECT 135.875 84.850 136.915 85.020 ;
        RECT 135.875 84.410 136.915 84.580 ;
        RECT 137.130 84.550 137.300 84.880 ;
        RECT 137.640 84.010 137.930 85.420 ;
        RECT 134.980 83.890 137.930 84.010 ;
        RECT 153.600 85.420 156.470 85.520 ;
        RECT 153.600 84.010 153.900 85.420 ;
        RECT 154.240 84.550 154.410 84.880 ;
        RECT 154.580 84.850 155.620 85.020 ;
        RECT 154.580 84.410 155.620 84.580 ;
        RECT 155.790 84.550 155.960 84.880 ;
        RECT 156.300 84.010 156.470 85.420 ;
        RECT 134.980 83.840 137.810 83.890 ;
        RECT 153.600 83.870 156.470 84.010 ;
        RECT 153.730 83.840 156.470 83.870 ;
        RECT 157.030 85.550 159.860 85.600 ;
        RECT 157.030 85.430 159.980 85.550 ;
        RECT 157.030 84.020 157.200 85.430 ;
        RECT 157.540 84.560 157.710 84.890 ;
        RECT 157.925 84.860 158.965 85.030 ;
        RECT 157.925 84.420 158.965 84.590 ;
        RECT 159.180 84.560 159.350 84.890 ;
        RECT 159.690 84.020 159.980 85.430 ;
        RECT 157.030 83.900 159.980 84.020 ;
        RECT 157.030 83.850 159.860 83.900 ;
        RECT 131.680 83.410 134.420 83.480 ;
        RECT 131.550 83.310 134.420 83.410 ;
        RECT 131.550 81.900 131.850 83.310 ;
        RECT 132.190 82.440 132.360 82.770 ;
        RECT 132.530 82.740 133.570 82.910 ;
        RECT 132.530 82.300 133.570 82.470 ;
        RECT 133.740 82.440 133.910 82.770 ;
        RECT 134.250 81.900 134.420 83.310 ;
        RECT 131.550 81.760 134.420 81.900 ;
        RECT 131.680 81.730 134.420 81.760 ;
        RECT 134.980 83.440 137.810 83.490 ;
        RECT 134.980 83.320 137.930 83.440 ;
        RECT 153.730 83.420 156.470 83.490 ;
        RECT 134.980 81.910 135.150 83.320 ;
        RECT 135.490 82.450 135.660 82.780 ;
        RECT 135.875 82.750 136.915 82.920 ;
        RECT 135.875 82.310 136.915 82.480 ;
        RECT 137.130 82.450 137.300 82.780 ;
        RECT 137.640 81.910 137.930 83.320 ;
        RECT 134.980 81.790 137.930 81.910 ;
        RECT 153.600 83.320 156.470 83.420 ;
        RECT 153.600 81.910 153.900 83.320 ;
        RECT 154.240 82.450 154.410 82.780 ;
        RECT 154.580 82.750 155.620 82.920 ;
        RECT 154.580 82.310 155.620 82.480 ;
        RECT 155.790 82.450 155.960 82.780 ;
        RECT 156.300 81.910 156.470 83.320 ;
        RECT 134.980 81.740 137.810 81.790 ;
        RECT 153.600 81.770 156.470 81.910 ;
        RECT 153.730 81.740 156.470 81.770 ;
        RECT 157.030 83.450 159.860 83.500 ;
        RECT 157.030 83.330 159.980 83.450 ;
        RECT 157.030 81.920 157.200 83.330 ;
        RECT 157.540 82.460 157.710 82.790 ;
        RECT 157.925 82.760 158.965 82.930 ;
        RECT 157.925 82.320 158.965 82.490 ;
        RECT 159.180 82.460 159.350 82.790 ;
        RECT 159.690 81.920 159.980 83.330 ;
        RECT 157.030 81.800 159.980 81.920 ;
        RECT 157.030 81.750 159.860 81.800 ;
        RECT 131.680 81.310 134.420 81.380 ;
        RECT 131.550 81.210 134.420 81.310 ;
        RECT 131.550 79.800 131.850 81.210 ;
        RECT 132.190 80.340 132.360 80.670 ;
        RECT 132.530 80.640 133.570 80.810 ;
        RECT 132.530 80.200 133.570 80.370 ;
        RECT 133.740 80.340 133.910 80.670 ;
        RECT 134.250 79.800 134.420 81.210 ;
        RECT 131.550 79.660 134.420 79.800 ;
        RECT 131.680 79.630 134.420 79.660 ;
        RECT 134.980 81.340 137.810 81.390 ;
        RECT 134.980 81.220 137.930 81.340 ;
        RECT 153.730 81.320 156.470 81.390 ;
        RECT 134.980 79.810 135.150 81.220 ;
        RECT 135.490 80.350 135.660 80.680 ;
        RECT 135.875 80.650 136.915 80.820 ;
        RECT 135.875 80.210 136.915 80.380 ;
        RECT 137.130 80.350 137.300 80.680 ;
        RECT 137.640 79.810 137.930 81.220 ;
        RECT 134.980 79.690 137.930 79.810 ;
        RECT 153.600 81.220 156.470 81.320 ;
        RECT 153.600 79.810 153.900 81.220 ;
        RECT 154.240 80.350 154.410 80.680 ;
        RECT 154.580 80.650 155.620 80.820 ;
        RECT 154.580 80.210 155.620 80.380 ;
        RECT 155.790 80.350 155.960 80.680 ;
        RECT 156.300 79.810 156.470 81.220 ;
        RECT 134.980 79.640 137.810 79.690 ;
        RECT 153.600 79.670 156.470 79.810 ;
        RECT 153.730 79.640 156.470 79.670 ;
        RECT 157.030 81.350 159.860 81.400 ;
        RECT 157.030 81.230 159.980 81.350 ;
        RECT 157.030 79.820 157.200 81.230 ;
        RECT 157.540 80.360 157.710 80.690 ;
        RECT 157.925 80.660 158.965 80.830 ;
        RECT 157.925 80.220 158.965 80.390 ;
        RECT 159.180 80.360 159.350 80.690 ;
        RECT 159.690 79.820 159.980 81.230 ;
        RECT 157.030 79.700 159.980 79.820 ;
        RECT 157.030 79.650 159.860 79.700 ;
        RECT 131.680 79.210 134.420 79.280 ;
        RECT 131.550 79.110 134.420 79.210 ;
        RECT 131.550 77.700 131.850 79.110 ;
        RECT 132.190 78.240 132.360 78.570 ;
        RECT 132.530 78.540 133.570 78.710 ;
        RECT 132.530 78.100 133.570 78.270 ;
        RECT 133.740 78.240 133.910 78.570 ;
        RECT 134.250 77.700 134.420 79.110 ;
        RECT 131.550 77.560 134.420 77.700 ;
        RECT 131.680 77.530 134.420 77.560 ;
        RECT 134.980 79.240 137.810 79.290 ;
        RECT 134.980 79.120 137.930 79.240 ;
        RECT 153.730 79.220 156.470 79.290 ;
        RECT 134.980 77.710 135.150 79.120 ;
        RECT 135.490 78.250 135.660 78.580 ;
        RECT 135.875 78.550 136.915 78.720 ;
        RECT 135.875 78.110 136.915 78.280 ;
        RECT 137.130 78.250 137.300 78.580 ;
        RECT 137.640 77.710 137.930 79.120 ;
        RECT 134.980 77.590 137.930 77.710 ;
        RECT 153.600 79.120 156.470 79.220 ;
        RECT 153.600 77.710 153.900 79.120 ;
        RECT 154.240 78.250 154.410 78.580 ;
        RECT 154.580 78.550 155.620 78.720 ;
        RECT 154.580 78.110 155.620 78.280 ;
        RECT 155.790 78.250 155.960 78.580 ;
        RECT 156.300 77.710 156.470 79.120 ;
        RECT 134.980 77.540 137.810 77.590 ;
        RECT 153.600 77.570 156.470 77.710 ;
        RECT 153.730 77.540 156.470 77.570 ;
        RECT 157.030 79.250 159.860 79.300 ;
        RECT 157.030 79.130 159.980 79.250 ;
        RECT 157.030 77.720 157.200 79.130 ;
        RECT 157.540 78.260 157.710 78.590 ;
        RECT 157.925 78.560 158.965 78.730 ;
        RECT 157.925 78.120 158.965 78.290 ;
        RECT 159.180 78.260 159.350 78.590 ;
        RECT 159.690 77.720 159.980 79.130 ;
        RECT 157.030 77.600 159.980 77.720 ;
        RECT 157.030 77.550 159.860 77.600 ;
        RECT 131.680 77.110 134.420 77.180 ;
        RECT 131.550 77.010 134.420 77.110 ;
        RECT 131.550 75.600 131.850 77.010 ;
        RECT 132.190 76.140 132.360 76.470 ;
        RECT 132.530 76.440 133.570 76.610 ;
        RECT 132.530 76.000 133.570 76.170 ;
        RECT 133.740 76.140 133.910 76.470 ;
        RECT 134.250 75.600 134.420 77.010 ;
        RECT 131.550 75.460 134.420 75.600 ;
        RECT 131.680 75.430 134.420 75.460 ;
        RECT 134.980 77.140 137.810 77.190 ;
        RECT 134.980 77.020 137.930 77.140 ;
        RECT 153.730 77.120 156.470 77.190 ;
        RECT 134.980 75.610 135.150 77.020 ;
        RECT 135.490 76.150 135.660 76.480 ;
        RECT 135.875 76.450 136.915 76.620 ;
        RECT 135.875 76.010 136.915 76.180 ;
        RECT 137.130 76.150 137.300 76.480 ;
        RECT 137.640 75.610 137.930 77.020 ;
        RECT 134.980 75.490 137.930 75.610 ;
        RECT 153.600 77.020 156.470 77.120 ;
        RECT 153.600 75.610 153.900 77.020 ;
        RECT 154.240 76.150 154.410 76.480 ;
        RECT 154.580 76.450 155.620 76.620 ;
        RECT 154.580 76.010 155.620 76.180 ;
        RECT 155.790 76.150 155.960 76.480 ;
        RECT 156.300 75.610 156.470 77.020 ;
        RECT 134.980 75.440 137.810 75.490 ;
        RECT 153.600 75.470 156.470 75.610 ;
        RECT 153.730 75.440 156.470 75.470 ;
        RECT 157.030 77.150 159.860 77.200 ;
        RECT 157.030 77.030 159.980 77.150 ;
        RECT 157.030 75.620 157.200 77.030 ;
        RECT 157.540 76.160 157.710 76.490 ;
        RECT 157.925 76.460 158.965 76.630 ;
        RECT 157.925 76.020 158.965 76.190 ;
        RECT 159.180 76.160 159.350 76.490 ;
        RECT 159.690 75.620 159.980 77.030 ;
        RECT 157.030 75.500 159.980 75.620 ;
        RECT 157.030 75.450 159.860 75.500 ;
        RECT 131.680 75.010 134.420 75.080 ;
        RECT 131.550 74.910 134.420 75.010 ;
        RECT 131.550 73.500 131.850 74.910 ;
        RECT 132.190 74.040 132.360 74.370 ;
        RECT 132.530 74.340 133.570 74.510 ;
        RECT 132.530 73.900 133.570 74.070 ;
        RECT 133.740 74.040 133.910 74.370 ;
        RECT 134.250 73.500 134.420 74.910 ;
        RECT 131.550 73.360 134.420 73.500 ;
        RECT 131.680 73.330 134.420 73.360 ;
        RECT 134.980 75.040 137.810 75.090 ;
        RECT 134.980 74.920 137.930 75.040 ;
        RECT 153.730 75.020 156.470 75.090 ;
        RECT 134.980 73.510 135.150 74.920 ;
        RECT 135.490 74.050 135.660 74.380 ;
        RECT 135.875 74.350 136.915 74.520 ;
        RECT 135.875 73.910 136.915 74.080 ;
        RECT 137.130 74.050 137.300 74.380 ;
        RECT 137.640 73.510 137.930 74.920 ;
        RECT 134.980 73.390 137.930 73.510 ;
        RECT 153.600 74.920 156.470 75.020 ;
        RECT 153.600 73.510 153.900 74.920 ;
        RECT 154.240 74.050 154.410 74.380 ;
        RECT 154.580 74.350 155.620 74.520 ;
        RECT 154.580 73.910 155.620 74.080 ;
        RECT 155.790 74.050 155.960 74.380 ;
        RECT 156.300 73.510 156.470 74.920 ;
        RECT 134.980 73.340 137.810 73.390 ;
        RECT 153.600 73.370 156.470 73.510 ;
        RECT 153.730 73.340 156.470 73.370 ;
        RECT 157.030 75.050 159.860 75.100 ;
        RECT 157.030 74.930 159.980 75.050 ;
        RECT 157.030 73.520 157.200 74.930 ;
        RECT 157.540 74.060 157.710 74.390 ;
        RECT 157.925 74.360 158.965 74.530 ;
        RECT 157.925 73.920 158.965 74.090 ;
        RECT 159.180 74.060 159.350 74.390 ;
        RECT 159.690 73.520 159.980 74.930 ;
        RECT 157.030 73.400 159.980 73.520 ;
        RECT 157.030 73.350 159.860 73.400 ;
        RECT 131.680 72.910 134.420 72.980 ;
        RECT 131.550 72.810 134.420 72.910 ;
        RECT 131.550 71.400 131.850 72.810 ;
        RECT 132.190 71.940 132.360 72.270 ;
        RECT 132.530 72.240 133.570 72.410 ;
        RECT 132.530 71.800 133.570 71.970 ;
        RECT 133.740 71.940 133.910 72.270 ;
        RECT 134.250 71.400 134.420 72.810 ;
        RECT 131.550 71.260 134.420 71.400 ;
        RECT 131.680 71.230 134.420 71.260 ;
        RECT 134.980 72.940 137.810 72.990 ;
        RECT 134.980 72.820 137.930 72.940 ;
        RECT 153.730 72.920 156.470 72.990 ;
        RECT 134.980 71.410 135.150 72.820 ;
        RECT 135.490 71.950 135.660 72.280 ;
        RECT 135.875 72.250 136.915 72.420 ;
        RECT 135.875 71.810 136.915 71.980 ;
        RECT 137.130 71.950 137.300 72.280 ;
        RECT 137.640 71.410 137.930 72.820 ;
        RECT 134.980 71.290 137.930 71.410 ;
        RECT 153.600 72.820 156.470 72.920 ;
        RECT 153.600 71.410 153.900 72.820 ;
        RECT 154.240 71.950 154.410 72.280 ;
        RECT 154.580 72.250 155.620 72.420 ;
        RECT 154.580 71.810 155.620 71.980 ;
        RECT 155.790 71.950 155.960 72.280 ;
        RECT 156.300 71.410 156.470 72.820 ;
        RECT 134.980 71.240 137.810 71.290 ;
        RECT 153.600 71.270 156.470 71.410 ;
        RECT 153.730 71.240 156.470 71.270 ;
        RECT 157.030 72.950 159.860 73.000 ;
        RECT 157.030 72.830 159.980 72.950 ;
        RECT 157.030 71.420 157.200 72.830 ;
        RECT 157.540 71.960 157.710 72.290 ;
        RECT 157.925 72.260 158.965 72.430 ;
        RECT 157.925 71.820 158.965 71.990 ;
        RECT 159.180 71.960 159.350 72.290 ;
        RECT 159.690 71.420 159.980 72.830 ;
        RECT 157.030 71.300 159.980 71.420 ;
        RECT 157.030 71.250 159.860 71.300 ;
        RECT 131.680 70.810 134.420 70.880 ;
        RECT 131.550 70.710 134.420 70.810 ;
        RECT 131.550 69.300 131.850 70.710 ;
        RECT 132.190 69.840 132.360 70.170 ;
        RECT 132.530 70.140 133.570 70.310 ;
        RECT 132.530 69.700 133.570 69.870 ;
        RECT 133.740 69.840 133.910 70.170 ;
        RECT 134.250 69.300 134.420 70.710 ;
        RECT 131.550 69.160 134.420 69.300 ;
        RECT 131.680 69.130 134.420 69.160 ;
        RECT 134.980 70.840 137.810 70.890 ;
        RECT 134.980 70.720 137.930 70.840 ;
        RECT 153.730 70.820 156.470 70.890 ;
        RECT 134.980 69.310 135.150 70.720 ;
        RECT 135.490 69.850 135.660 70.180 ;
        RECT 135.875 70.150 136.915 70.320 ;
        RECT 135.875 69.710 136.915 69.880 ;
        RECT 137.130 69.850 137.300 70.180 ;
        RECT 137.640 69.310 137.930 70.720 ;
        RECT 134.980 69.190 137.930 69.310 ;
        RECT 153.600 70.720 156.470 70.820 ;
        RECT 153.600 69.310 153.900 70.720 ;
        RECT 154.240 69.850 154.410 70.180 ;
        RECT 154.580 70.150 155.620 70.320 ;
        RECT 154.580 69.710 155.620 69.880 ;
        RECT 155.790 69.850 155.960 70.180 ;
        RECT 156.300 69.310 156.470 70.720 ;
        RECT 134.980 69.140 137.810 69.190 ;
        RECT 153.600 69.170 156.470 69.310 ;
        RECT 153.730 69.140 156.470 69.170 ;
        RECT 157.030 70.850 159.860 70.900 ;
        RECT 157.030 70.730 159.980 70.850 ;
        RECT 157.030 69.320 157.200 70.730 ;
        RECT 157.540 69.860 157.710 70.190 ;
        RECT 157.925 70.160 158.965 70.330 ;
        RECT 157.925 69.720 158.965 69.890 ;
        RECT 159.180 69.860 159.350 70.190 ;
        RECT 159.690 69.320 159.980 70.730 ;
        RECT 157.030 69.200 159.980 69.320 ;
        RECT 157.030 69.150 159.860 69.200 ;
        RECT 131.680 68.710 134.420 68.780 ;
        RECT 131.550 68.610 134.420 68.710 ;
        RECT 131.550 67.200 131.850 68.610 ;
        RECT 132.190 67.740 132.360 68.070 ;
        RECT 132.530 68.040 133.570 68.210 ;
        RECT 132.530 67.600 133.570 67.770 ;
        RECT 133.740 67.740 133.910 68.070 ;
        RECT 134.250 67.200 134.420 68.610 ;
        RECT 131.550 67.060 134.420 67.200 ;
        RECT 131.680 67.030 134.420 67.060 ;
        RECT 134.980 68.740 137.810 68.790 ;
        RECT 134.980 68.620 137.930 68.740 ;
        RECT 153.730 68.720 156.470 68.790 ;
        RECT 134.980 67.210 135.150 68.620 ;
        RECT 135.490 67.750 135.660 68.080 ;
        RECT 135.875 68.050 136.915 68.220 ;
        RECT 135.875 67.610 136.915 67.780 ;
        RECT 137.130 67.750 137.300 68.080 ;
        RECT 137.640 67.210 137.930 68.620 ;
        RECT 134.980 67.090 137.930 67.210 ;
        RECT 153.600 68.620 156.470 68.720 ;
        RECT 153.600 67.210 153.900 68.620 ;
        RECT 154.240 67.750 154.410 68.080 ;
        RECT 154.580 68.050 155.620 68.220 ;
        RECT 154.580 67.610 155.620 67.780 ;
        RECT 155.790 67.750 155.960 68.080 ;
        RECT 156.300 67.210 156.470 68.620 ;
        RECT 134.980 67.040 137.810 67.090 ;
        RECT 153.600 67.070 156.470 67.210 ;
        RECT 153.730 67.040 156.470 67.070 ;
        RECT 157.030 68.750 159.860 68.800 ;
        RECT 157.030 68.630 159.980 68.750 ;
        RECT 157.030 67.220 157.200 68.630 ;
        RECT 157.540 67.760 157.710 68.090 ;
        RECT 157.925 68.060 158.965 68.230 ;
        RECT 157.925 67.620 158.965 67.790 ;
        RECT 159.180 67.760 159.350 68.090 ;
        RECT 159.690 67.220 159.980 68.630 ;
        RECT 157.030 67.100 159.980 67.220 ;
        RECT 157.030 67.050 159.860 67.100 ;
        RECT 131.680 66.610 134.420 66.680 ;
        RECT 131.550 66.510 134.420 66.610 ;
        RECT 131.550 65.100 131.850 66.510 ;
        RECT 132.190 65.640 132.360 65.970 ;
        RECT 132.530 65.940 133.570 66.110 ;
        RECT 132.530 65.500 133.570 65.670 ;
        RECT 133.740 65.640 133.910 65.970 ;
        RECT 134.250 65.100 134.420 66.510 ;
        RECT 131.550 64.960 134.420 65.100 ;
        RECT 131.680 64.930 134.420 64.960 ;
        RECT 134.980 66.640 137.810 66.690 ;
        RECT 134.980 66.520 137.930 66.640 ;
        RECT 153.730 66.620 156.470 66.690 ;
        RECT 134.980 65.110 135.150 66.520 ;
        RECT 135.490 65.650 135.660 65.980 ;
        RECT 135.875 65.950 136.915 66.120 ;
        RECT 135.875 65.510 136.915 65.680 ;
        RECT 137.130 65.650 137.300 65.980 ;
        RECT 137.640 65.110 137.930 66.520 ;
        RECT 134.980 64.990 137.930 65.110 ;
        RECT 153.600 66.520 156.470 66.620 ;
        RECT 153.600 65.110 153.900 66.520 ;
        RECT 154.240 65.650 154.410 65.980 ;
        RECT 154.580 65.950 155.620 66.120 ;
        RECT 154.580 65.510 155.620 65.680 ;
        RECT 155.790 65.650 155.960 65.980 ;
        RECT 156.300 65.110 156.470 66.520 ;
        RECT 134.980 64.940 137.810 64.990 ;
        RECT 153.600 64.970 156.470 65.110 ;
        RECT 153.730 64.940 156.470 64.970 ;
        RECT 157.030 66.650 159.860 66.700 ;
        RECT 157.030 66.530 159.980 66.650 ;
        RECT 157.030 65.120 157.200 66.530 ;
        RECT 157.540 65.660 157.710 65.990 ;
        RECT 157.925 65.960 158.965 66.130 ;
        RECT 157.925 65.520 158.965 65.690 ;
        RECT 159.180 65.660 159.350 65.990 ;
        RECT 159.690 65.120 159.980 66.530 ;
        RECT 157.030 65.000 159.980 65.120 ;
        RECT 157.030 64.950 159.860 65.000 ;
        RECT 131.680 64.510 134.420 64.580 ;
        RECT 131.550 64.410 134.420 64.510 ;
        RECT 131.550 63.000 131.850 64.410 ;
        RECT 132.190 63.540 132.360 63.870 ;
        RECT 132.530 63.840 133.570 64.010 ;
        RECT 132.530 63.400 133.570 63.570 ;
        RECT 133.740 63.540 133.910 63.870 ;
        RECT 134.250 63.000 134.420 64.410 ;
        RECT 131.550 62.860 134.420 63.000 ;
        RECT 131.680 62.830 134.420 62.860 ;
        RECT 134.980 64.540 137.810 64.590 ;
        RECT 134.980 64.420 137.930 64.540 ;
        RECT 153.730 64.520 156.470 64.590 ;
        RECT 134.980 63.010 135.150 64.420 ;
        RECT 135.490 63.550 135.660 63.880 ;
        RECT 135.875 63.850 136.915 64.020 ;
        RECT 135.875 63.410 136.915 63.580 ;
        RECT 137.130 63.550 137.300 63.880 ;
        RECT 137.640 63.010 137.930 64.420 ;
        RECT 134.980 62.890 137.930 63.010 ;
        RECT 153.600 64.420 156.470 64.520 ;
        RECT 153.600 63.010 153.900 64.420 ;
        RECT 154.240 63.550 154.410 63.880 ;
        RECT 154.580 63.850 155.620 64.020 ;
        RECT 154.580 63.410 155.620 63.580 ;
        RECT 155.790 63.550 155.960 63.880 ;
        RECT 156.300 63.010 156.470 64.420 ;
        RECT 134.980 62.840 137.810 62.890 ;
        RECT 153.600 62.870 156.470 63.010 ;
        RECT 153.730 62.840 156.470 62.870 ;
        RECT 157.030 64.550 159.860 64.600 ;
        RECT 157.030 64.430 159.980 64.550 ;
        RECT 157.030 63.020 157.200 64.430 ;
        RECT 157.540 63.560 157.710 63.890 ;
        RECT 157.925 63.860 158.965 64.030 ;
        RECT 157.925 63.420 158.965 63.590 ;
        RECT 159.180 63.560 159.350 63.890 ;
        RECT 159.690 63.020 159.980 64.430 ;
        RECT 157.030 62.900 159.980 63.020 ;
        RECT 157.030 62.850 159.860 62.900 ;
        RECT 131.680 62.410 134.420 62.480 ;
        RECT 131.550 62.310 134.420 62.410 ;
        RECT 131.550 60.900 131.850 62.310 ;
        RECT 132.190 61.440 132.360 61.770 ;
        RECT 132.530 61.740 133.570 61.910 ;
        RECT 132.530 61.300 133.570 61.470 ;
        RECT 133.740 61.440 133.910 61.770 ;
        RECT 134.250 60.900 134.420 62.310 ;
        RECT 131.550 60.760 134.420 60.900 ;
        RECT 131.680 60.730 134.420 60.760 ;
        RECT 134.980 62.440 137.810 62.490 ;
        RECT 134.980 62.320 137.930 62.440 ;
        RECT 153.730 62.420 156.470 62.490 ;
        RECT 134.980 60.910 135.150 62.320 ;
        RECT 135.490 61.450 135.660 61.780 ;
        RECT 135.875 61.750 136.915 61.920 ;
        RECT 135.875 61.310 136.915 61.480 ;
        RECT 137.130 61.450 137.300 61.780 ;
        RECT 137.640 60.910 137.930 62.320 ;
        RECT 134.980 60.790 137.930 60.910 ;
        RECT 153.600 62.320 156.470 62.420 ;
        RECT 153.600 60.910 153.900 62.320 ;
        RECT 154.240 61.450 154.410 61.780 ;
        RECT 154.580 61.750 155.620 61.920 ;
        RECT 154.580 61.310 155.620 61.480 ;
        RECT 155.790 61.450 155.960 61.780 ;
        RECT 156.300 60.910 156.470 62.320 ;
        RECT 134.980 60.740 137.810 60.790 ;
        RECT 153.600 60.770 156.470 60.910 ;
        RECT 153.730 60.740 156.470 60.770 ;
        RECT 157.030 62.450 159.860 62.500 ;
        RECT 157.030 62.330 159.980 62.450 ;
        RECT 157.030 60.920 157.200 62.330 ;
        RECT 157.540 61.460 157.710 61.790 ;
        RECT 157.925 61.760 158.965 61.930 ;
        RECT 157.925 61.320 158.965 61.490 ;
        RECT 159.180 61.460 159.350 61.790 ;
        RECT 159.690 60.920 159.980 62.330 ;
        RECT 157.030 60.800 159.980 60.920 ;
        RECT 157.030 60.750 159.860 60.800 ;
        RECT 131.680 60.310 134.420 60.380 ;
        RECT 131.550 60.210 134.420 60.310 ;
        RECT 131.550 58.800 131.850 60.210 ;
        RECT 132.190 59.340 132.360 59.670 ;
        RECT 132.530 59.640 133.570 59.810 ;
        RECT 132.530 59.200 133.570 59.370 ;
        RECT 133.740 59.340 133.910 59.670 ;
        RECT 134.250 58.800 134.420 60.210 ;
        RECT 131.550 58.660 134.420 58.800 ;
        RECT 131.680 58.630 134.420 58.660 ;
        RECT 134.980 60.340 137.810 60.390 ;
        RECT 134.980 60.220 137.930 60.340 ;
        RECT 153.730 60.320 156.470 60.390 ;
        RECT 134.980 58.810 135.150 60.220 ;
        RECT 135.490 59.350 135.660 59.680 ;
        RECT 135.875 59.650 136.915 59.820 ;
        RECT 135.875 59.210 136.915 59.380 ;
        RECT 137.130 59.350 137.300 59.680 ;
        RECT 137.640 58.810 137.930 60.220 ;
        RECT 134.980 58.690 137.930 58.810 ;
        RECT 153.600 60.220 156.470 60.320 ;
        RECT 153.600 58.810 153.900 60.220 ;
        RECT 154.240 59.350 154.410 59.680 ;
        RECT 154.580 59.650 155.620 59.820 ;
        RECT 154.580 59.210 155.620 59.380 ;
        RECT 155.790 59.350 155.960 59.680 ;
        RECT 156.300 58.810 156.470 60.220 ;
        RECT 134.980 58.640 137.810 58.690 ;
        RECT 153.600 58.670 156.470 58.810 ;
        RECT 153.730 58.640 156.470 58.670 ;
        RECT 157.030 60.350 159.860 60.400 ;
        RECT 157.030 60.230 159.980 60.350 ;
        RECT 157.030 58.820 157.200 60.230 ;
        RECT 157.540 59.360 157.710 59.690 ;
        RECT 157.925 59.660 158.965 59.830 ;
        RECT 157.925 59.220 158.965 59.390 ;
        RECT 159.180 59.360 159.350 59.690 ;
        RECT 159.690 58.820 159.980 60.230 ;
        RECT 157.030 58.700 159.980 58.820 ;
        RECT 157.030 58.650 159.860 58.700 ;
        RECT 131.680 58.210 134.420 58.280 ;
        RECT 131.550 58.110 134.420 58.210 ;
        RECT 131.550 56.700 131.850 58.110 ;
        RECT 132.190 57.240 132.360 57.570 ;
        RECT 132.530 57.540 133.570 57.710 ;
        RECT 132.530 57.100 133.570 57.270 ;
        RECT 133.740 57.240 133.910 57.570 ;
        RECT 134.250 56.700 134.420 58.110 ;
        RECT 131.550 56.560 134.420 56.700 ;
        RECT 131.680 56.530 134.420 56.560 ;
        RECT 134.980 58.240 137.810 58.290 ;
        RECT 134.980 58.120 137.930 58.240 ;
        RECT 153.730 58.220 156.470 58.290 ;
        RECT 134.980 56.710 135.150 58.120 ;
        RECT 135.490 57.250 135.660 57.580 ;
        RECT 135.875 57.550 136.915 57.720 ;
        RECT 135.875 57.110 136.915 57.280 ;
        RECT 137.130 57.250 137.300 57.580 ;
        RECT 137.640 56.710 137.930 58.120 ;
        RECT 134.980 56.590 137.930 56.710 ;
        RECT 153.600 58.120 156.470 58.220 ;
        RECT 153.600 56.710 153.900 58.120 ;
        RECT 154.240 57.250 154.410 57.580 ;
        RECT 154.580 57.550 155.620 57.720 ;
        RECT 154.580 57.110 155.620 57.280 ;
        RECT 155.790 57.250 155.960 57.580 ;
        RECT 156.300 56.710 156.470 58.120 ;
        RECT 134.980 56.540 137.810 56.590 ;
        RECT 153.600 56.570 156.470 56.710 ;
        RECT 153.730 56.540 156.470 56.570 ;
        RECT 157.030 58.250 159.860 58.300 ;
        RECT 157.030 58.130 159.980 58.250 ;
        RECT 157.030 56.720 157.200 58.130 ;
        RECT 157.540 57.260 157.710 57.590 ;
        RECT 157.925 57.560 158.965 57.730 ;
        RECT 157.925 57.120 158.965 57.290 ;
        RECT 159.180 57.260 159.350 57.590 ;
        RECT 159.690 56.720 159.980 58.130 ;
        RECT 157.030 56.600 159.980 56.720 ;
        RECT 157.030 56.550 159.860 56.600 ;
        RECT 131.680 56.110 134.420 56.180 ;
        RECT 131.550 56.010 134.420 56.110 ;
        RECT 131.550 54.600 131.850 56.010 ;
        RECT 132.190 55.140 132.360 55.470 ;
        RECT 132.530 55.440 133.570 55.610 ;
        RECT 132.530 55.000 133.570 55.170 ;
        RECT 133.740 55.140 133.910 55.470 ;
        RECT 134.250 54.600 134.420 56.010 ;
        RECT 131.550 54.460 134.420 54.600 ;
        RECT 131.680 54.430 134.420 54.460 ;
        RECT 134.980 56.140 137.810 56.190 ;
        RECT 134.980 56.020 137.930 56.140 ;
        RECT 153.730 56.120 156.470 56.190 ;
        RECT 134.980 54.610 135.150 56.020 ;
        RECT 135.490 55.150 135.660 55.480 ;
        RECT 135.875 55.450 136.915 55.620 ;
        RECT 135.875 55.010 136.915 55.180 ;
        RECT 137.130 55.150 137.300 55.480 ;
        RECT 137.640 54.610 137.930 56.020 ;
        RECT 134.980 54.490 137.930 54.610 ;
        RECT 153.600 56.020 156.470 56.120 ;
        RECT 153.600 54.610 153.900 56.020 ;
        RECT 154.240 55.150 154.410 55.480 ;
        RECT 154.580 55.450 155.620 55.620 ;
        RECT 154.580 55.010 155.620 55.180 ;
        RECT 155.790 55.150 155.960 55.480 ;
        RECT 156.300 54.610 156.470 56.020 ;
        RECT 134.980 54.440 137.810 54.490 ;
        RECT 153.600 54.470 156.470 54.610 ;
        RECT 153.730 54.440 156.470 54.470 ;
        RECT 157.030 56.150 159.860 56.200 ;
        RECT 157.030 56.030 159.980 56.150 ;
        RECT 157.030 54.620 157.200 56.030 ;
        RECT 157.540 55.160 157.710 55.490 ;
        RECT 157.925 55.460 158.965 55.630 ;
        RECT 157.925 55.020 158.965 55.190 ;
        RECT 159.180 55.160 159.350 55.490 ;
        RECT 159.690 54.620 159.980 56.030 ;
        RECT 157.030 54.500 159.980 54.620 ;
        RECT 157.030 54.450 159.860 54.500 ;
        RECT 131.680 54.010 134.420 54.080 ;
        RECT 131.550 53.910 134.420 54.010 ;
        RECT 131.550 52.500 131.850 53.910 ;
        RECT 132.190 53.040 132.360 53.370 ;
        RECT 132.530 53.340 133.570 53.510 ;
        RECT 132.530 52.900 133.570 53.070 ;
        RECT 133.740 53.040 133.910 53.370 ;
        RECT 134.250 52.500 134.420 53.910 ;
        RECT 131.550 52.360 134.420 52.500 ;
        RECT 131.680 52.330 134.420 52.360 ;
        RECT 134.980 54.040 137.810 54.090 ;
        RECT 134.980 53.920 137.930 54.040 ;
        RECT 153.730 54.020 156.470 54.090 ;
        RECT 134.980 52.510 135.150 53.920 ;
        RECT 135.490 53.050 135.660 53.380 ;
        RECT 135.875 53.350 136.915 53.520 ;
        RECT 135.875 52.910 136.915 53.080 ;
        RECT 137.130 53.050 137.300 53.380 ;
        RECT 137.640 52.510 137.930 53.920 ;
        RECT 134.980 52.390 137.930 52.510 ;
        RECT 153.600 53.920 156.470 54.020 ;
        RECT 153.600 52.510 153.900 53.920 ;
        RECT 154.240 53.050 154.410 53.380 ;
        RECT 154.580 53.350 155.620 53.520 ;
        RECT 154.580 52.910 155.620 53.080 ;
        RECT 155.790 53.050 155.960 53.380 ;
        RECT 156.300 52.510 156.470 53.920 ;
        RECT 134.980 52.340 137.810 52.390 ;
        RECT 153.600 52.370 156.470 52.510 ;
        RECT 153.730 52.340 156.470 52.370 ;
        RECT 157.030 54.050 159.860 54.100 ;
        RECT 157.030 53.930 159.980 54.050 ;
        RECT 157.030 52.520 157.200 53.930 ;
        RECT 157.540 53.060 157.710 53.390 ;
        RECT 157.925 53.360 158.965 53.530 ;
        RECT 157.925 52.920 158.965 53.090 ;
        RECT 159.180 53.060 159.350 53.390 ;
        RECT 159.690 52.520 159.980 53.930 ;
        RECT 157.030 52.400 159.980 52.520 ;
        RECT 157.030 52.350 159.860 52.400 ;
        RECT 131.680 51.910 134.420 51.980 ;
        RECT 131.550 51.810 134.420 51.910 ;
        RECT 131.550 50.400 131.850 51.810 ;
        RECT 132.190 50.940 132.360 51.270 ;
        RECT 132.530 51.240 133.570 51.410 ;
        RECT 132.530 50.800 133.570 50.970 ;
        RECT 133.740 50.940 133.910 51.270 ;
        RECT 134.250 50.400 134.420 51.810 ;
        RECT 131.550 50.260 134.420 50.400 ;
        RECT 131.680 50.230 134.420 50.260 ;
        RECT 134.980 51.940 137.810 51.990 ;
        RECT 134.980 51.820 137.930 51.940 ;
        RECT 153.730 51.920 156.470 51.990 ;
        RECT 134.980 50.410 135.150 51.820 ;
        RECT 135.490 50.950 135.660 51.280 ;
        RECT 135.875 51.250 136.915 51.420 ;
        RECT 135.875 50.810 136.915 50.980 ;
        RECT 137.130 50.950 137.300 51.280 ;
        RECT 137.640 50.410 137.930 51.820 ;
        RECT 134.980 50.290 137.930 50.410 ;
        RECT 153.600 51.820 156.470 51.920 ;
        RECT 153.600 50.410 153.900 51.820 ;
        RECT 154.240 50.950 154.410 51.280 ;
        RECT 154.580 51.250 155.620 51.420 ;
        RECT 154.580 50.810 155.620 50.980 ;
        RECT 155.790 50.950 155.960 51.280 ;
        RECT 156.300 50.410 156.470 51.820 ;
        RECT 134.980 50.240 137.810 50.290 ;
        RECT 153.600 50.270 156.470 50.410 ;
        RECT 153.730 50.240 156.470 50.270 ;
        RECT 157.030 51.950 159.860 52.000 ;
        RECT 157.030 51.830 159.980 51.950 ;
        RECT 157.030 50.420 157.200 51.830 ;
        RECT 157.540 50.960 157.710 51.290 ;
        RECT 157.925 51.260 158.965 51.430 ;
        RECT 157.925 50.820 158.965 50.990 ;
        RECT 159.180 50.960 159.350 51.290 ;
        RECT 159.690 50.420 159.980 51.830 ;
        RECT 157.030 50.300 159.980 50.420 ;
        RECT 157.030 50.250 159.860 50.300 ;
        RECT 131.680 49.810 134.420 49.880 ;
        RECT 131.550 49.710 134.420 49.810 ;
        RECT 131.550 48.300 131.850 49.710 ;
        RECT 132.190 48.840 132.360 49.170 ;
        RECT 132.530 49.140 133.570 49.310 ;
        RECT 132.530 48.700 133.570 48.870 ;
        RECT 133.740 48.840 133.910 49.170 ;
        RECT 134.250 48.300 134.420 49.710 ;
        RECT 131.550 48.160 134.420 48.300 ;
        RECT 131.680 48.130 134.420 48.160 ;
        RECT 134.980 49.840 137.810 49.890 ;
        RECT 134.980 49.720 137.930 49.840 ;
        RECT 153.730 49.820 156.470 49.890 ;
        RECT 134.980 48.310 135.150 49.720 ;
        RECT 135.490 48.850 135.660 49.180 ;
        RECT 135.875 49.150 136.915 49.320 ;
        RECT 135.875 48.710 136.915 48.880 ;
        RECT 137.130 48.850 137.300 49.180 ;
        RECT 137.640 48.310 137.930 49.720 ;
        RECT 134.980 48.190 137.930 48.310 ;
        RECT 153.600 49.720 156.470 49.820 ;
        RECT 153.600 48.310 153.900 49.720 ;
        RECT 154.240 48.850 154.410 49.180 ;
        RECT 154.580 49.150 155.620 49.320 ;
        RECT 154.580 48.710 155.620 48.880 ;
        RECT 155.790 48.850 155.960 49.180 ;
        RECT 156.300 48.310 156.470 49.720 ;
        RECT 134.980 48.140 137.810 48.190 ;
        RECT 153.600 48.170 156.470 48.310 ;
        RECT 153.730 48.140 156.470 48.170 ;
        RECT 157.030 49.850 159.860 49.900 ;
        RECT 157.030 49.730 159.980 49.850 ;
        RECT 157.030 48.320 157.200 49.730 ;
        RECT 157.540 48.860 157.710 49.190 ;
        RECT 157.925 49.160 158.965 49.330 ;
        RECT 157.925 48.720 158.965 48.890 ;
        RECT 159.180 48.860 159.350 49.190 ;
        RECT 159.690 48.320 159.980 49.730 ;
        RECT 157.030 48.200 159.980 48.320 ;
        RECT 157.030 48.150 159.860 48.200 ;
        RECT 131.680 47.710 134.420 47.780 ;
        RECT 131.550 47.610 134.420 47.710 ;
        RECT 131.550 46.200 131.850 47.610 ;
        RECT 132.190 46.740 132.360 47.070 ;
        RECT 132.530 47.040 133.570 47.210 ;
        RECT 132.530 46.600 133.570 46.770 ;
        RECT 133.740 46.740 133.910 47.070 ;
        RECT 134.250 46.200 134.420 47.610 ;
        RECT 131.550 46.060 134.420 46.200 ;
        RECT 131.680 46.030 134.420 46.060 ;
        RECT 134.980 47.740 137.810 47.790 ;
        RECT 134.980 47.620 137.930 47.740 ;
        RECT 153.730 47.720 156.470 47.790 ;
        RECT 134.980 46.210 135.150 47.620 ;
        RECT 135.490 46.750 135.660 47.080 ;
        RECT 135.875 47.050 136.915 47.220 ;
        RECT 135.875 46.610 136.915 46.780 ;
        RECT 137.130 46.750 137.300 47.080 ;
        RECT 137.640 46.210 137.930 47.620 ;
        RECT 134.980 46.090 137.930 46.210 ;
        RECT 153.600 47.620 156.470 47.720 ;
        RECT 153.600 46.210 153.900 47.620 ;
        RECT 154.240 46.750 154.410 47.080 ;
        RECT 154.580 47.050 155.620 47.220 ;
        RECT 154.580 46.610 155.620 46.780 ;
        RECT 155.790 46.750 155.960 47.080 ;
        RECT 156.300 46.210 156.470 47.620 ;
        RECT 134.980 46.040 137.810 46.090 ;
        RECT 153.600 46.070 156.470 46.210 ;
        RECT 153.730 46.040 156.470 46.070 ;
        RECT 157.030 47.750 159.860 47.800 ;
        RECT 157.030 47.630 159.980 47.750 ;
        RECT 157.030 46.220 157.200 47.630 ;
        RECT 157.540 46.760 157.710 47.090 ;
        RECT 157.925 47.060 158.965 47.230 ;
        RECT 157.925 46.620 158.965 46.790 ;
        RECT 159.180 46.760 159.350 47.090 ;
        RECT 159.690 46.220 159.980 47.630 ;
        RECT 157.030 46.100 159.980 46.220 ;
        RECT 157.030 46.050 159.860 46.100 ;
        RECT 131.680 45.610 134.420 45.680 ;
        RECT 131.550 45.510 134.420 45.610 ;
        RECT 131.550 44.100 131.850 45.510 ;
        RECT 132.190 44.640 132.360 44.970 ;
        RECT 132.530 44.940 133.570 45.110 ;
        RECT 132.530 44.500 133.570 44.670 ;
        RECT 133.740 44.640 133.910 44.970 ;
        RECT 134.250 44.100 134.420 45.510 ;
        RECT 131.550 43.960 134.420 44.100 ;
        RECT 131.680 43.930 134.420 43.960 ;
        RECT 134.980 45.640 137.810 45.690 ;
        RECT 134.980 45.520 137.930 45.640 ;
        RECT 153.730 45.620 156.470 45.690 ;
        RECT 134.980 44.110 135.150 45.520 ;
        RECT 135.490 44.650 135.660 44.980 ;
        RECT 135.875 44.950 136.915 45.120 ;
        RECT 135.875 44.510 136.915 44.680 ;
        RECT 137.130 44.650 137.300 44.980 ;
        RECT 137.640 44.110 137.930 45.520 ;
        RECT 134.980 43.990 137.930 44.110 ;
        RECT 153.600 45.520 156.470 45.620 ;
        RECT 153.600 44.110 153.900 45.520 ;
        RECT 154.240 44.650 154.410 44.980 ;
        RECT 154.580 44.950 155.620 45.120 ;
        RECT 154.580 44.510 155.620 44.680 ;
        RECT 155.790 44.650 155.960 44.980 ;
        RECT 156.300 44.110 156.470 45.520 ;
        RECT 134.980 43.940 137.810 43.990 ;
        RECT 153.600 43.970 156.470 44.110 ;
        RECT 153.730 43.940 156.470 43.970 ;
        RECT 157.030 45.650 159.860 45.700 ;
        RECT 157.030 45.530 159.980 45.650 ;
        RECT 157.030 44.120 157.200 45.530 ;
        RECT 157.540 44.660 157.710 44.990 ;
        RECT 157.925 44.960 158.965 45.130 ;
        RECT 157.925 44.520 158.965 44.690 ;
        RECT 159.180 44.660 159.350 44.990 ;
        RECT 159.690 44.120 159.980 45.530 ;
        RECT 157.030 44.000 159.980 44.120 ;
        RECT 157.030 43.950 159.860 44.000 ;
        RECT 131.680 43.510 134.420 43.580 ;
        RECT 131.550 43.410 134.420 43.510 ;
        RECT 131.550 42.000 131.850 43.410 ;
        RECT 132.190 42.540 132.360 42.870 ;
        RECT 132.530 42.840 133.570 43.010 ;
        RECT 132.530 42.400 133.570 42.570 ;
        RECT 133.740 42.540 133.910 42.870 ;
        RECT 134.250 42.000 134.420 43.410 ;
        RECT 131.550 41.860 134.420 42.000 ;
        RECT 131.680 41.830 134.420 41.860 ;
        RECT 134.980 43.540 137.810 43.590 ;
        RECT 134.980 43.420 137.930 43.540 ;
        RECT 153.730 43.520 156.470 43.590 ;
        RECT 134.980 42.010 135.150 43.420 ;
        RECT 135.490 42.550 135.660 42.880 ;
        RECT 135.875 42.850 136.915 43.020 ;
        RECT 135.875 42.410 136.915 42.580 ;
        RECT 137.130 42.550 137.300 42.880 ;
        RECT 137.640 42.010 137.930 43.420 ;
        RECT 134.980 41.890 137.930 42.010 ;
        RECT 153.600 43.420 156.470 43.520 ;
        RECT 153.600 42.010 153.900 43.420 ;
        RECT 154.240 42.550 154.410 42.880 ;
        RECT 154.580 42.850 155.620 43.020 ;
        RECT 154.580 42.410 155.620 42.580 ;
        RECT 155.790 42.550 155.960 42.880 ;
        RECT 156.300 42.010 156.470 43.420 ;
        RECT 134.980 41.840 137.810 41.890 ;
        RECT 153.600 41.870 156.470 42.010 ;
        RECT 153.730 41.840 156.470 41.870 ;
        RECT 157.030 43.550 159.860 43.600 ;
        RECT 157.030 43.430 159.980 43.550 ;
        RECT 157.030 42.020 157.200 43.430 ;
        RECT 157.540 42.560 157.710 42.890 ;
        RECT 157.925 42.860 158.965 43.030 ;
        RECT 157.925 42.420 158.965 42.590 ;
        RECT 159.180 42.560 159.350 42.890 ;
        RECT 159.690 42.020 159.980 43.430 ;
        RECT 157.030 41.900 159.980 42.020 ;
        RECT 157.030 41.850 159.860 41.900 ;
        RECT 131.680 41.410 134.420 41.480 ;
        RECT 131.550 41.310 134.420 41.410 ;
        RECT 131.550 39.900 131.850 41.310 ;
        RECT 132.190 40.440 132.360 40.770 ;
        RECT 132.530 40.740 133.570 40.910 ;
        RECT 132.530 40.300 133.570 40.470 ;
        RECT 133.740 40.440 133.910 40.770 ;
        RECT 134.250 39.900 134.420 41.310 ;
        RECT 131.550 39.760 134.420 39.900 ;
        RECT 131.680 39.730 134.420 39.760 ;
        RECT 134.980 41.440 137.810 41.490 ;
        RECT 134.980 41.320 137.930 41.440 ;
        RECT 153.730 41.420 156.470 41.490 ;
        RECT 134.980 39.910 135.150 41.320 ;
        RECT 135.490 40.450 135.660 40.780 ;
        RECT 135.875 40.750 136.915 40.920 ;
        RECT 135.875 40.310 136.915 40.480 ;
        RECT 137.130 40.450 137.300 40.780 ;
        RECT 137.640 39.910 137.930 41.320 ;
        RECT 134.980 39.790 137.930 39.910 ;
        RECT 153.600 41.320 156.470 41.420 ;
        RECT 153.600 39.910 153.900 41.320 ;
        RECT 154.240 40.450 154.410 40.780 ;
        RECT 154.580 40.750 155.620 40.920 ;
        RECT 154.580 40.310 155.620 40.480 ;
        RECT 155.790 40.450 155.960 40.780 ;
        RECT 156.300 39.910 156.470 41.320 ;
        RECT 134.980 39.740 137.810 39.790 ;
        RECT 153.600 39.770 156.470 39.910 ;
        RECT 153.730 39.740 156.470 39.770 ;
        RECT 157.030 41.450 159.860 41.500 ;
        RECT 157.030 41.330 159.980 41.450 ;
        RECT 157.030 39.920 157.200 41.330 ;
        RECT 157.540 40.460 157.710 40.790 ;
        RECT 157.925 40.760 158.965 40.930 ;
        RECT 157.925 40.320 158.965 40.490 ;
        RECT 159.180 40.460 159.350 40.790 ;
        RECT 159.690 39.920 159.980 41.330 ;
        RECT 157.030 39.800 159.980 39.920 ;
        RECT 157.030 39.750 159.860 39.800 ;
        RECT 131.680 39.310 134.420 39.380 ;
        RECT 131.550 39.210 134.420 39.310 ;
        RECT 131.550 37.800 131.850 39.210 ;
        RECT 132.190 38.340 132.360 38.670 ;
        RECT 132.530 38.640 133.570 38.810 ;
        RECT 132.530 38.200 133.570 38.370 ;
        RECT 133.740 38.340 133.910 38.670 ;
        RECT 134.250 37.800 134.420 39.210 ;
        RECT 131.550 37.660 134.420 37.800 ;
        RECT 131.680 37.630 134.420 37.660 ;
        RECT 134.980 39.340 137.810 39.390 ;
        RECT 134.980 39.220 137.930 39.340 ;
        RECT 153.730 39.320 156.470 39.390 ;
        RECT 134.980 37.810 135.150 39.220 ;
        RECT 135.490 38.350 135.660 38.680 ;
        RECT 135.875 38.650 136.915 38.820 ;
        RECT 135.875 38.210 136.915 38.380 ;
        RECT 137.130 38.350 137.300 38.680 ;
        RECT 137.640 37.810 137.930 39.220 ;
        RECT 134.980 37.690 137.930 37.810 ;
        RECT 153.600 39.220 156.470 39.320 ;
        RECT 153.600 37.810 153.900 39.220 ;
        RECT 154.240 38.350 154.410 38.680 ;
        RECT 154.580 38.650 155.620 38.820 ;
        RECT 154.580 38.210 155.620 38.380 ;
        RECT 155.790 38.350 155.960 38.680 ;
        RECT 156.300 37.810 156.470 39.220 ;
        RECT 134.980 37.640 137.810 37.690 ;
        RECT 153.600 37.670 156.470 37.810 ;
        RECT 153.730 37.640 156.470 37.670 ;
        RECT 157.030 39.350 159.860 39.400 ;
        RECT 157.030 39.230 159.980 39.350 ;
        RECT 157.030 37.820 157.200 39.230 ;
        RECT 157.540 38.360 157.710 38.690 ;
        RECT 157.925 38.660 158.965 38.830 ;
        RECT 157.925 38.220 158.965 38.390 ;
        RECT 159.180 38.360 159.350 38.690 ;
        RECT 159.690 37.820 159.980 39.230 ;
        RECT 157.030 37.700 159.980 37.820 ;
        RECT 157.030 37.650 159.860 37.700 ;
        RECT 131.680 37.210 134.420 37.280 ;
        RECT 131.550 37.110 134.420 37.210 ;
        RECT 131.550 35.700 131.850 37.110 ;
        RECT 132.190 36.240 132.360 36.570 ;
        RECT 132.530 36.540 133.570 36.710 ;
        RECT 132.530 36.100 133.570 36.270 ;
        RECT 133.740 36.240 133.910 36.570 ;
        RECT 134.250 35.700 134.420 37.110 ;
        RECT 131.550 35.560 134.420 35.700 ;
        RECT 131.680 35.530 134.420 35.560 ;
        RECT 134.980 37.240 137.810 37.290 ;
        RECT 134.980 37.120 137.930 37.240 ;
        RECT 153.730 37.220 156.470 37.290 ;
        RECT 134.980 35.710 135.150 37.120 ;
        RECT 135.490 36.250 135.660 36.580 ;
        RECT 135.875 36.550 136.915 36.720 ;
        RECT 135.875 36.110 136.915 36.280 ;
        RECT 137.130 36.250 137.300 36.580 ;
        RECT 137.640 35.710 137.930 37.120 ;
        RECT 134.980 35.590 137.930 35.710 ;
        RECT 153.600 37.120 156.470 37.220 ;
        RECT 153.600 35.710 153.900 37.120 ;
        RECT 154.240 36.250 154.410 36.580 ;
        RECT 154.580 36.550 155.620 36.720 ;
        RECT 154.580 36.110 155.620 36.280 ;
        RECT 155.790 36.250 155.960 36.580 ;
        RECT 156.300 35.710 156.470 37.120 ;
        RECT 134.980 35.540 137.810 35.590 ;
        RECT 153.600 35.570 156.470 35.710 ;
        RECT 153.730 35.540 156.470 35.570 ;
        RECT 157.030 37.250 159.860 37.300 ;
        RECT 157.030 37.130 159.980 37.250 ;
        RECT 157.030 35.720 157.200 37.130 ;
        RECT 157.540 36.260 157.710 36.590 ;
        RECT 157.925 36.560 158.965 36.730 ;
        RECT 157.925 36.120 158.965 36.290 ;
        RECT 159.180 36.260 159.350 36.590 ;
        RECT 159.690 35.720 159.980 37.130 ;
        RECT 157.030 35.600 159.980 35.720 ;
        RECT 157.030 35.550 159.860 35.600 ;
        RECT 131.680 35.110 134.420 35.180 ;
        RECT 131.550 35.010 134.420 35.110 ;
        RECT 131.550 33.600 131.850 35.010 ;
        RECT 132.190 34.140 132.360 34.470 ;
        RECT 132.530 34.440 133.570 34.610 ;
        RECT 132.530 34.000 133.570 34.170 ;
        RECT 133.740 34.140 133.910 34.470 ;
        RECT 134.250 33.600 134.420 35.010 ;
        RECT 131.550 33.460 134.420 33.600 ;
        RECT 131.680 33.430 134.420 33.460 ;
        RECT 134.980 35.140 137.810 35.190 ;
        RECT 134.980 35.020 137.930 35.140 ;
        RECT 153.730 35.120 156.470 35.190 ;
        RECT 134.980 33.610 135.150 35.020 ;
        RECT 135.490 34.150 135.660 34.480 ;
        RECT 135.875 34.450 136.915 34.620 ;
        RECT 135.875 34.010 136.915 34.180 ;
        RECT 137.130 34.150 137.300 34.480 ;
        RECT 137.640 33.610 137.930 35.020 ;
        RECT 134.980 33.490 137.930 33.610 ;
        RECT 153.600 35.020 156.470 35.120 ;
        RECT 153.600 33.610 153.900 35.020 ;
        RECT 154.240 34.150 154.410 34.480 ;
        RECT 154.580 34.450 155.620 34.620 ;
        RECT 154.580 34.010 155.620 34.180 ;
        RECT 155.790 34.150 155.960 34.480 ;
        RECT 156.300 33.610 156.470 35.020 ;
        RECT 134.980 33.440 137.810 33.490 ;
        RECT 153.600 33.470 156.470 33.610 ;
        RECT 153.730 33.440 156.470 33.470 ;
        RECT 157.030 35.150 159.860 35.200 ;
        RECT 157.030 35.030 159.980 35.150 ;
        RECT 157.030 33.620 157.200 35.030 ;
        RECT 157.540 34.160 157.710 34.490 ;
        RECT 157.925 34.460 158.965 34.630 ;
        RECT 157.925 34.020 158.965 34.190 ;
        RECT 159.180 34.160 159.350 34.490 ;
        RECT 159.690 33.620 159.980 35.030 ;
        RECT 157.030 33.500 159.980 33.620 ;
        RECT 157.030 33.450 159.860 33.500 ;
        RECT 131.680 33.010 134.420 33.080 ;
        RECT 131.550 32.910 134.420 33.010 ;
        RECT 131.550 31.500 131.850 32.910 ;
        RECT 132.190 32.040 132.360 32.370 ;
        RECT 132.530 32.340 133.570 32.510 ;
        RECT 132.530 31.900 133.570 32.070 ;
        RECT 133.740 32.040 133.910 32.370 ;
        RECT 134.250 31.500 134.420 32.910 ;
        RECT 131.550 31.360 134.420 31.500 ;
        RECT 131.680 31.330 134.420 31.360 ;
        RECT 134.980 33.040 137.810 33.090 ;
        RECT 134.980 32.920 137.930 33.040 ;
        RECT 153.730 33.020 156.470 33.090 ;
        RECT 134.980 31.510 135.150 32.920 ;
        RECT 135.490 32.050 135.660 32.380 ;
        RECT 135.875 32.350 136.915 32.520 ;
        RECT 135.875 31.910 136.915 32.080 ;
        RECT 137.130 32.050 137.300 32.380 ;
        RECT 137.640 31.510 137.930 32.920 ;
        RECT 134.980 31.390 137.930 31.510 ;
        RECT 153.600 32.920 156.470 33.020 ;
        RECT 153.600 31.510 153.900 32.920 ;
        RECT 154.240 32.050 154.410 32.380 ;
        RECT 154.580 32.350 155.620 32.520 ;
        RECT 154.580 31.910 155.620 32.080 ;
        RECT 155.790 32.050 155.960 32.380 ;
        RECT 156.300 31.510 156.470 32.920 ;
        RECT 134.980 31.340 137.810 31.390 ;
        RECT 153.600 31.370 156.470 31.510 ;
        RECT 153.730 31.340 156.470 31.370 ;
        RECT 157.030 33.050 159.860 33.100 ;
        RECT 157.030 32.930 159.980 33.050 ;
        RECT 157.030 31.520 157.200 32.930 ;
        RECT 157.540 32.060 157.710 32.390 ;
        RECT 157.925 32.360 158.965 32.530 ;
        RECT 157.925 31.920 158.965 32.090 ;
        RECT 159.180 32.060 159.350 32.390 ;
        RECT 159.690 31.520 159.980 32.930 ;
        RECT 157.030 31.400 159.980 31.520 ;
        RECT 157.030 31.350 159.860 31.400 ;
        RECT 131.680 30.910 134.420 30.980 ;
        RECT 131.550 30.810 134.420 30.910 ;
        RECT 131.550 29.400 131.850 30.810 ;
        RECT 132.190 29.940 132.360 30.270 ;
        RECT 132.530 30.240 133.570 30.410 ;
        RECT 132.530 29.800 133.570 29.970 ;
        RECT 133.740 29.940 133.910 30.270 ;
        RECT 134.250 29.400 134.420 30.810 ;
        RECT 131.550 29.260 134.420 29.400 ;
        RECT 131.680 29.230 134.420 29.260 ;
        RECT 134.980 30.940 137.810 30.990 ;
        RECT 134.980 30.820 137.930 30.940 ;
        RECT 153.730 30.920 156.470 30.990 ;
        RECT 134.980 29.410 135.150 30.820 ;
        RECT 135.490 29.950 135.660 30.280 ;
        RECT 135.875 30.250 136.915 30.420 ;
        RECT 135.875 29.810 136.915 29.980 ;
        RECT 137.130 29.950 137.300 30.280 ;
        RECT 137.640 29.410 137.930 30.820 ;
        RECT 134.980 29.290 137.930 29.410 ;
        RECT 153.600 30.820 156.470 30.920 ;
        RECT 153.600 29.410 153.900 30.820 ;
        RECT 154.240 29.950 154.410 30.280 ;
        RECT 154.580 30.250 155.620 30.420 ;
        RECT 154.580 29.810 155.620 29.980 ;
        RECT 155.790 29.950 155.960 30.280 ;
        RECT 156.300 29.410 156.470 30.820 ;
        RECT 134.980 29.240 137.810 29.290 ;
        RECT 153.600 29.270 156.470 29.410 ;
        RECT 153.730 29.240 156.470 29.270 ;
        RECT 157.030 30.950 159.860 31.000 ;
        RECT 157.030 30.830 159.980 30.950 ;
        RECT 157.030 29.420 157.200 30.830 ;
        RECT 157.540 29.960 157.710 30.290 ;
        RECT 157.925 30.260 158.965 30.430 ;
        RECT 157.925 29.820 158.965 29.990 ;
        RECT 159.180 29.960 159.350 30.290 ;
        RECT 159.690 29.420 159.980 30.830 ;
        RECT 157.030 29.300 159.980 29.420 ;
        RECT 157.030 29.250 159.860 29.300 ;
        RECT 131.680 28.810 134.420 28.880 ;
        RECT 131.550 28.710 134.420 28.810 ;
        RECT 131.550 27.300 131.850 28.710 ;
        RECT 132.190 27.840 132.360 28.170 ;
        RECT 132.530 28.140 133.570 28.310 ;
        RECT 132.530 27.700 133.570 27.870 ;
        RECT 133.740 27.840 133.910 28.170 ;
        RECT 134.250 27.300 134.420 28.710 ;
        RECT 131.550 27.160 134.420 27.300 ;
        RECT 131.680 27.130 134.420 27.160 ;
        RECT 134.980 28.840 137.810 28.890 ;
        RECT 134.980 28.720 137.930 28.840 ;
        RECT 153.730 28.820 156.470 28.890 ;
        RECT 134.980 27.310 135.150 28.720 ;
        RECT 135.490 27.850 135.660 28.180 ;
        RECT 135.875 28.150 136.915 28.320 ;
        RECT 135.875 27.710 136.915 27.880 ;
        RECT 137.130 27.850 137.300 28.180 ;
        RECT 137.640 27.310 137.930 28.720 ;
        RECT 134.980 27.190 137.930 27.310 ;
        RECT 153.600 28.720 156.470 28.820 ;
        RECT 153.600 27.310 153.900 28.720 ;
        RECT 154.240 27.850 154.410 28.180 ;
        RECT 154.580 28.150 155.620 28.320 ;
        RECT 154.580 27.710 155.620 27.880 ;
        RECT 155.790 27.850 155.960 28.180 ;
        RECT 156.300 27.310 156.470 28.720 ;
        RECT 134.980 27.140 137.810 27.190 ;
        RECT 153.600 27.170 156.470 27.310 ;
        RECT 153.730 27.140 156.470 27.170 ;
        RECT 157.030 28.850 159.860 28.900 ;
        RECT 157.030 28.730 159.980 28.850 ;
        RECT 157.030 27.320 157.200 28.730 ;
        RECT 157.540 27.860 157.710 28.190 ;
        RECT 157.925 28.160 158.965 28.330 ;
        RECT 157.925 27.720 158.965 27.890 ;
        RECT 159.180 27.860 159.350 28.190 ;
        RECT 159.690 27.320 159.980 28.730 ;
        RECT 157.030 27.200 159.980 27.320 ;
        RECT 157.030 27.150 159.860 27.200 ;
        RECT 131.680 26.710 134.420 26.780 ;
        RECT 131.550 26.610 134.420 26.710 ;
        RECT 131.550 25.200 131.850 26.610 ;
        RECT 132.190 25.740 132.360 26.070 ;
        RECT 132.530 26.040 133.570 26.210 ;
        RECT 132.530 25.600 133.570 25.770 ;
        RECT 133.740 25.740 133.910 26.070 ;
        RECT 134.250 25.200 134.420 26.610 ;
        RECT 131.550 25.060 134.420 25.200 ;
        RECT 131.680 25.030 134.420 25.060 ;
        RECT 134.980 26.740 137.810 26.790 ;
        RECT 134.980 26.620 137.930 26.740 ;
        RECT 153.730 26.720 156.470 26.790 ;
        RECT 134.980 25.210 135.150 26.620 ;
        RECT 135.490 25.750 135.660 26.080 ;
        RECT 135.875 26.050 136.915 26.220 ;
        RECT 135.875 25.610 136.915 25.780 ;
        RECT 137.130 25.750 137.300 26.080 ;
        RECT 137.640 25.210 137.930 26.620 ;
        RECT 134.980 25.090 137.930 25.210 ;
        RECT 153.600 26.620 156.470 26.720 ;
        RECT 153.600 25.210 153.900 26.620 ;
        RECT 154.240 25.750 154.410 26.080 ;
        RECT 154.580 26.050 155.620 26.220 ;
        RECT 154.580 25.610 155.620 25.780 ;
        RECT 155.790 25.750 155.960 26.080 ;
        RECT 156.300 25.210 156.470 26.620 ;
        RECT 134.980 25.040 137.810 25.090 ;
        RECT 153.600 25.070 156.470 25.210 ;
        RECT 153.730 25.040 156.470 25.070 ;
        RECT 157.030 26.750 159.860 26.800 ;
        RECT 157.030 26.630 159.980 26.750 ;
        RECT 157.030 25.220 157.200 26.630 ;
        RECT 157.540 25.760 157.710 26.090 ;
        RECT 157.925 26.060 158.965 26.230 ;
        RECT 157.925 25.620 158.965 25.790 ;
        RECT 159.180 25.760 159.350 26.090 ;
        RECT 159.690 25.220 159.980 26.630 ;
        RECT 157.030 25.100 159.980 25.220 ;
        RECT 157.030 25.050 159.860 25.100 ;
        RECT 131.680 24.610 134.420 24.680 ;
        RECT 131.550 24.510 134.420 24.610 ;
        RECT 131.550 23.100 131.850 24.510 ;
        RECT 132.190 23.640 132.360 23.970 ;
        RECT 132.530 23.940 133.570 24.110 ;
        RECT 132.530 23.500 133.570 23.670 ;
        RECT 133.740 23.640 133.910 23.970 ;
        RECT 134.250 23.100 134.420 24.510 ;
        RECT 131.550 22.960 134.420 23.100 ;
        RECT 131.680 22.930 134.420 22.960 ;
        RECT 134.980 24.640 137.810 24.690 ;
        RECT 134.980 24.520 137.930 24.640 ;
        RECT 153.730 24.620 156.470 24.690 ;
        RECT 134.980 23.110 135.150 24.520 ;
        RECT 135.490 23.650 135.660 23.980 ;
        RECT 135.875 23.950 136.915 24.120 ;
        RECT 135.875 23.510 136.915 23.680 ;
        RECT 137.130 23.650 137.300 23.980 ;
        RECT 137.640 23.110 137.930 24.520 ;
        RECT 134.980 22.990 137.930 23.110 ;
        RECT 153.600 24.520 156.470 24.620 ;
        RECT 153.600 23.110 153.900 24.520 ;
        RECT 154.240 23.650 154.410 23.980 ;
        RECT 154.580 23.950 155.620 24.120 ;
        RECT 154.580 23.510 155.620 23.680 ;
        RECT 155.790 23.650 155.960 23.980 ;
        RECT 156.300 23.110 156.470 24.520 ;
        RECT 134.980 22.940 137.810 22.990 ;
        RECT 153.600 22.970 156.470 23.110 ;
        RECT 153.730 22.940 156.470 22.970 ;
        RECT 157.030 24.650 159.860 24.700 ;
        RECT 157.030 24.530 159.980 24.650 ;
        RECT 157.030 23.120 157.200 24.530 ;
        RECT 157.540 23.660 157.710 23.990 ;
        RECT 157.925 23.960 158.965 24.130 ;
        RECT 157.925 23.520 158.965 23.690 ;
        RECT 159.180 23.660 159.350 23.990 ;
        RECT 159.690 23.120 159.980 24.530 ;
        RECT 157.030 23.000 159.980 23.120 ;
        RECT 157.030 22.950 159.860 23.000 ;
        RECT 131.680 22.510 134.420 22.580 ;
        RECT 131.550 22.410 134.420 22.510 ;
        RECT 131.550 21.000 131.850 22.410 ;
        RECT 132.190 21.540 132.360 21.870 ;
        RECT 132.530 21.840 133.570 22.010 ;
        RECT 132.530 21.400 133.570 21.570 ;
        RECT 133.740 21.540 133.910 21.870 ;
        RECT 134.250 21.000 134.420 22.410 ;
        RECT 131.550 20.860 134.420 21.000 ;
        RECT 131.680 20.830 134.420 20.860 ;
        RECT 134.980 22.540 137.810 22.590 ;
        RECT 134.980 22.420 137.930 22.540 ;
        RECT 153.730 22.520 156.470 22.590 ;
        RECT 134.980 21.010 135.150 22.420 ;
        RECT 135.490 21.550 135.660 21.880 ;
        RECT 135.875 21.850 136.915 22.020 ;
        RECT 135.875 21.410 136.915 21.580 ;
        RECT 137.130 21.550 137.300 21.880 ;
        RECT 137.640 21.010 137.930 22.420 ;
        RECT 134.980 20.890 137.930 21.010 ;
        RECT 153.600 22.420 156.470 22.520 ;
        RECT 153.600 21.010 153.900 22.420 ;
        RECT 154.240 21.550 154.410 21.880 ;
        RECT 154.580 21.850 155.620 22.020 ;
        RECT 154.580 21.410 155.620 21.580 ;
        RECT 155.790 21.550 155.960 21.880 ;
        RECT 156.300 21.010 156.470 22.420 ;
        RECT 134.980 20.840 137.810 20.890 ;
        RECT 153.600 20.870 156.470 21.010 ;
        RECT 153.730 20.840 156.470 20.870 ;
        RECT 157.030 22.550 159.860 22.600 ;
        RECT 157.030 22.430 159.980 22.550 ;
        RECT 157.030 21.020 157.200 22.430 ;
        RECT 157.540 21.560 157.710 21.890 ;
        RECT 157.925 21.860 158.965 22.030 ;
        RECT 157.925 21.420 158.965 21.590 ;
        RECT 159.180 21.560 159.350 21.890 ;
        RECT 159.690 21.020 159.980 22.430 ;
        RECT 157.030 20.900 159.980 21.020 ;
        RECT 157.030 20.850 159.860 20.900 ;
        RECT 131.680 20.410 134.420 20.480 ;
        RECT 131.550 20.310 134.420 20.410 ;
        RECT 131.550 18.900 131.850 20.310 ;
        RECT 132.190 19.440 132.360 19.770 ;
        RECT 132.530 19.740 133.570 19.910 ;
        RECT 132.530 19.300 133.570 19.470 ;
        RECT 133.740 19.440 133.910 19.770 ;
        RECT 134.250 18.900 134.420 20.310 ;
        RECT 131.550 18.760 134.420 18.900 ;
        RECT 131.680 18.730 134.420 18.760 ;
        RECT 134.980 20.440 137.810 20.490 ;
        RECT 134.980 20.320 137.930 20.440 ;
        RECT 153.730 20.420 156.470 20.490 ;
        RECT 134.980 18.910 135.150 20.320 ;
        RECT 135.490 19.450 135.660 19.780 ;
        RECT 135.875 19.750 136.915 19.920 ;
        RECT 135.875 19.310 136.915 19.480 ;
        RECT 137.130 19.450 137.300 19.780 ;
        RECT 137.640 18.910 137.930 20.320 ;
        RECT 134.980 18.790 137.930 18.910 ;
        RECT 153.600 20.320 156.470 20.420 ;
        RECT 153.600 18.910 153.900 20.320 ;
        RECT 154.240 19.450 154.410 19.780 ;
        RECT 154.580 19.750 155.620 19.920 ;
        RECT 154.580 19.310 155.620 19.480 ;
        RECT 155.790 19.450 155.960 19.780 ;
        RECT 156.300 18.910 156.470 20.320 ;
        RECT 134.980 18.740 137.810 18.790 ;
        RECT 153.600 18.770 156.470 18.910 ;
        RECT 153.730 18.740 156.470 18.770 ;
        RECT 157.030 20.450 159.860 20.500 ;
        RECT 157.030 20.330 159.980 20.450 ;
        RECT 157.030 18.920 157.200 20.330 ;
        RECT 157.540 19.460 157.710 19.790 ;
        RECT 157.925 19.760 158.965 19.930 ;
        RECT 157.925 19.320 158.965 19.490 ;
        RECT 159.180 19.460 159.350 19.790 ;
        RECT 159.690 18.920 159.980 20.330 ;
        RECT 157.030 18.800 159.980 18.920 ;
        RECT 157.030 18.750 159.860 18.800 ;
        RECT 131.680 18.310 134.420 18.380 ;
        RECT 131.550 18.210 134.420 18.310 ;
        RECT 131.550 16.800 131.850 18.210 ;
        RECT 132.190 17.340 132.360 17.670 ;
        RECT 132.530 17.640 133.570 17.810 ;
        RECT 132.530 17.200 133.570 17.370 ;
        RECT 133.740 17.340 133.910 17.670 ;
        RECT 134.250 16.800 134.420 18.210 ;
        RECT 131.550 16.660 134.420 16.800 ;
        RECT 131.680 16.630 134.420 16.660 ;
        RECT 134.980 18.340 137.810 18.390 ;
        RECT 134.980 18.220 137.930 18.340 ;
        RECT 153.730 18.320 156.470 18.390 ;
        RECT 134.980 16.810 135.150 18.220 ;
        RECT 135.490 17.350 135.660 17.680 ;
        RECT 135.875 17.650 136.915 17.820 ;
        RECT 135.875 17.210 136.915 17.380 ;
        RECT 137.130 17.350 137.300 17.680 ;
        RECT 137.640 16.810 137.930 18.220 ;
        RECT 134.980 16.690 137.930 16.810 ;
        RECT 153.600 18.220 156.470 18.320 ;
        RECT 153.600 16.810 153.900 18.220 ;
        RECT 154.240 17.350 154.410 17.680 ;
        RECT 154.580 17.650 155.620 17.820 ;
        RECT 154.580 17.210 155.620 17.380 ;
        RECT 155.790 17.350 155.960 17.680 ;
        RECT 156.300 16.810 156.470 18.220 ;
        RECT 134.980 16.640 137.810 16.690 ;
        RECT 153.600 16.670 156.470 16.810 ;
        RECT 153.730 16.640 156.470 16.670 ;
        RECT 157.030 18.350 159.860 18.400 ;
        RECT 157.030 18.230 159.980 18.350 ;
        RECT 157.030 16.820 157.200 18.230 ;
        RECT 157.540 17.360 157.710 17.690 ;
        RECT 157.925 17.660 158.965 17.830 ;
        RECT 157.925 17.220 158.965 17.390 ;
        RECT 159.180 17.360 159.350 17.690 ;
        RECT 159.690 16.820 159.980 18.230 ;
        RECT 157.030 16.700 159.980 16.820 ;
        RECT 157.030 16.650 159.860 16.700 ;
        RECT 131.680 16.210 134.420 16.280 ;
        RECT 131.550 16.110 134.420 16.210 ;
        RECT 131.550 14.700 131.850 16.110 ;
        RECT 132.190 15.240 132.360 15.570 ;
        RECT 132.530 15.540 133.570 15.710 ;
        RECT 132.530 15.100 133.570 15.270 ;
        RECT 133.740 15.240 133.910 15.570 ;
        RECT 134.250 14.700 134.420 16.110 ;
        RECT 131.550 14.560 134.420 14.700 ;
        RECT 131.680 14.530 134.420 14.560 ;
        RECT 134.980 16.240 137.810 16.290 ;
        RECT 134.980 16.120 137.930 16.240 ;
        RECT 153.730 16.220 156.470 16.290 ;
        RECT 134.980 14.710 135.150 16.120 ;
        RECT 135.490 15.250 135.660 15.580 ;
        RECT 135.875 15.550 136.915 15.720 ;
        RECT 135.875 15.110 136.915 15.280 ;
        RECT 137.130 15.250 137.300 15.580 ;
        RECT 137.640 14.710 137.930 16.120 ;
        RECT 134.980 14.590 137.930 14.710 ;
        RECT 153.600 16.120 156.470 16.220 ;
        RECT 153.600 14.710 153.900 16.120 ;
        RECT 154.240 15.250 154.410 15.580 ;
        RECT 154.580 15.550 155.620 15.720 ;
        RECT 154.580 15.110 155.620 15.280 ;
        RECT 155.790 15.250 155.960 15.580 ;
        RECT 156.300 14.710 156.470 16.120 ;
        RECT 134.980 14.540 137.810 14.590 ;
        RECT 153.600 14.570 156.470 14.710 ;
        RECT 153.730 14.540 156.470 14.570 ;
        RECT 157.030 16.250 159.860 16.300 ;
        RECT 157.030 16.130 159.980 16.250 ;
        RECT 157.030 14.720 157.200 16.130 ;
        RECT 157.540 15.260 157.710 15.590 ;
        RECT 157.925 15.560 158.965 15.730 ;
        RECT 157.925 15.120 158.965 15.290 ;
        RECT 159.180 15.260 159.350 15.590 ;
        RECT 159.690 14.720 159.980 16.130 ;
        RECT 157.030 14.600 159.980 14.720 ;
        RECT 157.030 14.550 159.860 14.600 ;
        RECT 131.680 14.110 134.420 14.180 ;
        RECT 131.550 14.010 134.420 14.110 ;
        RECT 131.550 12.600 131.850 14.010 ;
        RECT 132.190 13.140 132.360 13.470 ;
        RECT 132.530 13.440 133.570 13.610 ;
        RECT 132.530 13.000 133.570 13.170 ;
        RECT 133.740 13.140 133.910 13.470 ;
        RECT 134.250 12.600 134.420 14.010 ;
        RECT 131.550 12.460 134.420 12.600 ;
        RECT 131.680 12.430 134.420 12.460 ;
        RECT 134.980 14.140 137.810 14.190 ;
        RECT 134.980 14.020 137.930 14.140 ;
        RECT 153.730 14.120 156.470 14.190 ;
        RECT 134.980 12.610 135.150 14.020 ;
        RECT 135.490 13.150 135.660 13.480 ;
        RECT 135.875 13.450 136.915 13.620 ;
        RECT 135.875 13.010 136.915 13.180 ;
        RECT 137.130 13.150 137.300 13.480 ;
        RECT 137.640 12.610 137.930 14.020 ;
        RECT 134.980 12.490 137.930 12.610 ;
        RECT 153.600 14.020 156.470 14.120 ;
        RECT 153.600 12.610 153.900 14.020 ;
        RECT 154.240 13.150 154.410 13.480 ;
        RECT 154.580 13.450 155.620 13.620 ;
        RECT 154.580 13.010 155.620 13.180 ;
        RECT 155.790 13.150 155.960 13.480 ;
        RECT 156.300 12.610 156.470 14.020 ;
        RECT 134.980 12.440 137.810 12.490 ;
        RECT 153.600 12.470 156.470 12.610 ;
        RECT 153.730 12.440 156.470 12.470 ;
        RECT 157.030 14.150 159.860 14.200 ;
        RECT 157.030 14.030 159.980 14.150 ;
        RECT 157.030 12.620 157.200 14.030 ;
        RECT 157.540 13.160 157.710 13.490 ;
        RECT 157.925 13.460 158.965 13.630 ;
        RECT 157.925 13.020 158.965 13.190 ;
        RECT 159.180 13.160 159.350 13.490 ;
        RECT 159.690 12.620 159.980 14.030 ;
        RECT 157.030 12.500 159.980 12.620 ;
        RECT 157.030 12.450 159.860 12.500 ;
        RECT 131.680 12.010 134.420 12.080 ;
        RECT 131.550 11.910 134.420 12.010 ;
        RECT 131.550 10.500 131.850 11.910 ;
        RECT 132.190 11.040 132.360 11.370 ;
        RECT 132.530 11.340 133.570 11.510 ;
        RECT 132.530 10.900 133.570 11.070 ;
        RECT 133.740 11.040 133.910 11.370 ;
        RECT 134.250 10.500 134.420 11.910 ;
        RECT 131.550 10.360 134.420 10.500 ;
        RECT 131.680 10.330 134.420 10.360 ;
        RECT 134.980 12.040 137.810 12.090 ;
        RECT 134.980 11.920 137.930 12.040 ;
        RECT 153.730 12.020 156.470 12.090 ;
        RECT 134.980 10.510 135.150 11.920 ;
        RECT 135.490 11.050 135.660 11.380 ;
        RECT 135.875 11.350 136.915 11.520 ;
        RECT 135.875 10.910 136.915 11.080 ;
        RECT 137.130 11.050 137.300 11.380 ;
        RECT 137.640 10.510 137.930 11.920 ;
        RECT 134.980 10.390 137.930 10.510 ;
        RECT 153.600 11.920 156.470 12.020 ;
        RECT 153.600 10.510 153.900 11.920 ;
        RECT 154.240 11.050 154.410 11.380 ;
        RECT 154.580 11.350 155.620 11.520 ;
        RECT 154.580 10.910 155.620 11.080 ;
        RECT 155.790 11.050 155.960 11.380 ;
        RECT 156.300 10.510 156.470 11.920 ;
        RECT 134.980 10.340 137.810 10.390 ;
        RECT 153.600 10.370 156.470 10.510 ;
        RECT 153.730 10.340 156.470 10.370 ;
        RECT 157.030 12.050 159.860 12.100 ;
        RECT 157.030 11.930 159.980 12.050 ;
        RECT 157.030 10.520 157.200 11.930 ;
        RECT 157.540 11.060 157.710 11.390 ;
        RECT 157.925 11.360 158.965 11.530 ;
        RECT 157.925 10.920 158.965 11.090 ;
        RECT 159.180 11.060 159.350 11.390 ;
        RECT 159.690 10.520 159.980 11.930 ;
        RECT 157.030 10.400 159.980 10.520 ;
        RECT 157.030 10.350 159.860 10.400 ;
        RECT 131.680 9.910 134.420 9.980 ;
        RECT 131.550 9.810 134.420 9.910 ;
        RECT 131.550 8.400 131.850 9.810 ;
        RECT 132.190 8.940 132.360 9.270 ;
        RECT 132.530 9.240 133.570 9.410 ;
        RECT 132.530 8.800 133.570 8.970 ;
        RECT 133.740 8.940 133.910 9.270 ;
        RECT 134.250 8.400 134.420 9.810 ;
        RECT 131.550 8.260 134.420 8.400 ;
        RECT 131.680 8.230 134.420 8.260 ;
        RECT 134.980 9.940 137.810 9.990 ;
        RECT 134.980 9.820 137.930 9.940 ;
        RECT 153.730 9.920 156.470 9.990 ;
        RECT 134.980 8.410 135.150 9.820 ;
        RECT 135.490 8.950 135.660 9.280 ;
        RECT 135.875 9.250 136.915 9.420 ;
        RECT 135.875 8.810 136.915 8.980 ;
        RECT 137.130 8.950 137.300 9.280 ;
        RECT 137.640 8.410 137.930 9.820 ;
        RECT 134.980 8.290 137.930 8.410 ;
        RECT 153.600 9.820 156.470 9.920 ;
        RECT 153.600 8.410 153.900 9.820 ;
        RECT 154.240 8.950 154.410 9.280 ;
        RECT 154.580 9.250 155.620 9.420 ;
        RECT 154.580 8.810 155.620 8.980 ;
        RECT 155.790 8.950 155.960 9.280 ;
        RECT 156.300 8.410 156.470 9.820 ;
        RECT 134.980 8.240 137.810 8.290 ;
        RECT 153.600 8.270 156.470 8.410 ;
        RECT 153.730 8.240 156.470 8.270 ;
        RECT 157.030 9.950 159.860 10.000 ;
        RECT 157.030 9.830 159.980 9.950 ;
        RECT 157.030 8.420 157.200 9.830 ;
        RECT 157.540 8.960 157.710 9.290 ;
        RECT 157.925 9.260 158.965 9.430 ;
        RECT 157.925 8.820 158.965 8.990 ;
        RECT 159.180 8.960 159.350 9.290 ;
        RECT 159.690 8.420 159.980 9.830 ;
        RECT 157.030 8.300 159.980 8.420 ;
        RECT 157.030 8.250 159.860 8.300 ;
        RECT 131.680 7.810 134.420 7.880 ;
        RECT 131.550 7.710 134.420 7.810 ;
        RECT 131.550 6.300 131.850 7.710 ;
        RECT 132.190 6.840 132.360 7.170 ;
        RECT 132.530 7.140 133.570 7.310 ;
        RECT 132.530 6.700 133.570 6.870 ;
        RECT 133.740 6.840 133.910 7.170 ;
        RECT 134.250 6.300 134.420 7.710 ;
        RECT 131.550 6.160 134.420 6.300 ;
        RECT 131.680 6.130 134.420 6.160 ;
        RECT 134.980 7.840 137.810 7.890 ;
        RECT 134.980 7.720 137.930 7.840 ;
        RECT 153.730 7.820 156.470 7.890 ;
        RECT 134.980 6.310 135.150 7.720 ;
        RECT 135.490 6.850 135.660 7.180 ;
        RECT 135.875 7.150 136.915 7.320 ;
        RECT 135.875 6.710 136.915 6.880 ;
        RECT 137.130 6.850 137.300 7.180 ;
        RECT 137.640 6.310 137.930 7.720 ;
        RECT 134.980 6.190 137.930 6.310 ;
        RECT 153.600 7.720 156.470 7.820 ;
        RECT 153.600 6.310 153.900 7.720 ;
        RECT 154.240 6.850 154.410 7.180 ;
        RECT 154.580 7.150 155.620 7.320 ;
        RECT 154.580 6.710 155.620 6.880 ;
        RECT 155.790 6.850 155.960 7.180 ;
        RECT 156.300 6.310 156.470 7.720 ;
        RECT 134.980 6.140 137.810 6.190 ;
        RECT 153.600 6.170 156.470 6.310 ;
        RECT 153.730 6.140 156.470 6.170 ;
        RECT 157.030 7.850 159.860 7.900 ;
        RECT 157.030 7.730 159.980 7.850 ;
        RECT 157.030 6.320 157.200 7.730 ;
        RECT 157.540 6.860 157.710 7.190 ;
        RECT 157.925 7.160 158.965 7.330 ;
        RECT 157.925 6.720 158.965 6.890 ;
        RECT 159.180 6.860 159.350 7.190 ;
        RECT 159.690 6.320 159.980 7.730 ;
        RECT 157.030 6.200 159.980 6.320 ;
        RECT 157.030 6.150 159.860 6.200 ;
        RECT 131.680 5.710 134.420 5.780 ;
        RECT 131.550 5.610 134.420 5.710 ;
        RECT 131.550 4.200 131.850 5.610 ;
        RECT 132.190 4.740 132.360 5.070 ;
        RECT 132.530 5.040 133.570 5.210 ;
        RECT 132.530 4.600 133.570 4.770 ;
        RECT 133.740 4.740 133.910 5.070 ;
        RECT 134.250 4.200 134.420 5.610 ;
        RECT 131.550 4.060 134.420 4.200 ;
        RECT 131.680 4.030 134.420 4.060 ;
        RECT 134.980 5.740 137.810 5.790 ;
        RECT 134.980 5.620 137.930 5.740 ;
        RECT 153.730 5.720 156.470 5.790 ;
        RECT 134.980 4.210 135.150 5.620 ;
        RECT 135.490 4.750 135.660 5.080 ;
        RECT 135.875 5.050 136.915 5.220 ;
        RECT 135.875 4.610 136.915 4.780 ;
        RECT 137.130 4.750 137.300 5.080 ;
        RECT 137.640 4.210 137.930 5.620 ;
        RECT 134.980 4.090 137.930 4.210 ;
        RECT 153.600 5.620 156.470 5.720 ;
        RECT 153.600 4.210 153.900 5.620 ;
        RECT 154.240 4.750 154.410 5.080 ;
        RECT 154.580 5.050 155.620 5.220 ;
        RECT 154.580 4.610 155.620 4.780 ;
        RECT 155.790 4.750 155.960 5.080 ;
        RECT 156.300 4.210 156.470 5.620 ;
        RECT 134.980 4.040 137.810 4.090 ;
        RECT 153.600 4.070 156.470 4.210 ;
        RECT 153.730 4.040 156.470 4.070 ;
        RECT 157.030 5.750 159.860 5.800 ;
        RECT 157.030 5.630 159.980 5.750 ;
        RECT 157.030 4.220 157.200 5.630 ;
        RECT 157.540 4.760 157.710 5.090 ;
        RECT 157.925 5.060 158.965 5.230 ;
        RECT 157.925 4.620 158.965 4.790 ;
        RECT 159.180 4.760 159.350 5.090 ;
        RECT 159.690 4.220 159.980 5.630 ;
        RECT 157.030 4.100 159.980 4.220 ;
        RECT 157.030 4.050 159.860 4.100 ;
        RECT 131.680 3.610 134.420 3.680 ;
        RECT 131.550 3.510 134.420 3.610 ;
        RECT 131.550 2.100 131.850 3.510 ;
        RECT 132.190 2.640 132.360 2.970 ;
        RECT 132.530 2.940 133.570 3.110 ;
        RECT 132.530 2.500 133.570 2.670 ;
        RECT 133.740 2.640 133.910 2.970 ;
        RECT 134.250 2.100 134.420 3.510 ;
        RECT 131.550 1.960 134.420 2.100 ;
        RECT 131.680 1.930 134.420 1.960 ;
        RECT 134.980 3.640 137.810 3.690 ;
        RECT 134.980 3.520 137.930 3.640 ;
        RECT 153.730 3.620 156.470 3.690 ;
        RECT 134.980 2.110 135.150 3.520 ;
        RECT 135.490 2.650 135.660 2.980 ;
        RECT 135.875 2.950 136.915 3.120 ;
        RECT 135.875 2.510 136.915 2.680 ;
        RECT 137.130 2.650 137.300 2.980 ;
        RECT 137.640 2.110 137.930 3.520 ;
        RECT 134.980 1.990 137.930 2.110 ;
        RECT 153.600 3.520 156.470 3.620 ;
        RECT 153.600 2.110 153.900 3.520 ;
        RECT 154.240 2.650 154.410 2.980 ;
        RECT 154.580 2.950 155.620 3.120 ;
        RECT 154.580 2.510 155.620 2.680 ;
        RECT 155.790 2.650 155.960 2.980 ;
        RECT 156.300 2.110 156.470 3.520 ;
        RECT 134.980 1.940 137.810 1.990 ;
        RECT 153.600 1.970 156.470 2.110 ;
        RECT 153.730 1.940 156.470 1.970 ;
        RECT 157.030 3.650 159.860 3.700 ;
        RECT 157.030 3.530 159.980 3.650 ;
        RECT 157.030 2.120 157.200 3.530 ;
        RECT 157.540 2.660 157.710 2.990 ;
        RECT 157.925 2.960 158.965 3.130 ;
        RECT 157.925 2.520 158.965 2.690 ;
        RECT 159.180 2.660 159.350 2.990 ;
        RECT 159.690 2.120 159.980 3.530 ;
        RECT 157.030 2.000 159.980 2.120 ;
        RECT 157.030 1.950 159.860 2.000 ;
      LAYER mcon ;
        RECT 132.610 210.780 133.490 210.950 ;
        RECT 132.190 210.560 132.360 210.730 ;
        RECT 133.740 210.560 133.910 210.730 ;
        RECT 132.610 210.340 133.490 210.510 ;
        RECT 135.955 210.790 136.835 210.960 ;
        RECT 135.490 210.570 135.660 210.740 ;
        RECT 137.130 210.570 137.300 210.740 ;
        RECT 135.955 210.350 136.835 210.520 ;
        RECT 137.670 209.830 137.930 211.480 ;
        RECT 154.660 210.850 155.540 211.020 ;
        RECT 154.240 210.630 154.410 210.800 ;
        RECT 155.790 210.630 155.960 210.800 ;
        RECT 154.660 210.410 155.540 210.580 ;
        RECT 158.005 210.860 158.885 211.030 ;
        RECT 157.540 210.640 157.710 210.810 ;
        RECT 159.180 210.640 159.350 210.810 ;
        RECT 158.005 210.420 158.885 210.590 ;
        RECT 159.720 209.900 159.980 211.550 ;
        RECT 132.610 208.680 133.490 208.850 ;
        RECT 132.190 208.460 132.360 208.630 ;
        RECT 133.740 208.460 133.910 208.630 ;
        RECT 132.610 208.240 133.490 208.410 ;
        RECT 135.955 208.690 136.835 208.860 ;
        RECT 135.490 208.470 135.660 208.640 ;
        RECT 137.130 208.470 137.300 208.640 ;
        RECT 135.955 208.250 136.835 208.420 ;
        RECT 137.670 207.730 137.930 209.380 ;
        RECT 154.660 208.750 155.540 208.920 ;
        RECT 154.240 208.530 154.410 208.700 ;
        RECT 155.790 208.530 155.960 208.700 ;
        RECT 154.660 208.310 155.540 208.480 ;
        RECT 158.005 208.760 158.885 208.930 ;
        RECT 157.540 208.540 157.710 208.710 ;
        RECT 159.180 208.540 159.350 208.710 ;
        RECT 158.005 208.320 158.885 208.490 ;
        RECT 159.720 207.800 159.980 209.450 ;
        RECT 132.610 206.580 133.490 206.750 ;
        RECT 132.190 206.360 132.360 206.530 ;
        RECT 133.740 206.360 133.910 206.530 ;
        RECT 132.610 206.140 133.490 206.310 ;
        RECT 135.955 206.590 136.835 206.760 ;
        RECT 135.490 206.370 135.660 206.540 ;
        RECT 137.130 206.370 137.300 206.540 ;
        RECT 135.955 206.150 136.835 206.320 ;
        RECT 137.670 205.630 137.930 207.280 ;
        RECT 154.660 206.650 155.540 206.820 ;
        RECT 154.240 206.430 154.410 206.600 ;
        RECT 155.790 206.430 155.960 206.600 ;
        RECT 154.660 206.210 155.540 206.380 ;
        RECT 158.005 206.660 158.885 206.830 ;
        RECT 157.540 206.440 157.710 206.610 ;
        RECT 159.180 206.440 159.350 206.610 ;
        RECT 158.005 206.220 158.885 206.390 ;
        RECT 159.720 205.700 159.980 207.350 ;
        RECT 132.610 204.480 133.490 204.650 ;
        RECT 132.190 204.260 132.360 204.430 ;
        RECT 133.740 204.260 133.910 204.430 ;
        RECT 132.610 204.040 133.490 204.210 ;
        RECT 135.955 204.490 136.835 204.660 ;
        RECT 135.490 204.270 135.660 204.440 ;
        RECT 137.130 204.270 137.300 204.440 ;
        RECT 135.955 204.050 136.835 204.220 ;
        RECT 137.670 203.530 137.930 205.180 ;
        RECT 154.660 204.550 155.540 204.720 ;
        RECT 154.240 204.330 154.410 204.500 ;
        RECT 155.790 204.330 155.960 204.500 ;
        RECT 154.660 204.110 155.540 204.280 ;
        RECT 158.005 204.560 158.885 204.730 ;
        RECT 157.540 204.340 157.710 204.510 ;
        RECT 159.180 204.340 159.350 204.510 ;
        RECT 158.005 204.120 158.885 204.290 ;
        RECT 159.720 203.600 159.980 205.250 ;
        RECT 132.610 202.390 133.490 202.560 ;
        RECT 132.190 202.170 132.360 202.340 ;
        RECT 133.740 202.170 133.910 202.340 ;
        RECT 132.610 201.950 133.490 202.120 ;
        RECT 135.955 202.400 136.835 202.570 ;
        RECT 135.490 202.180 135.660 202.350 ;
        RECT 137.130 202.180 137.300 202.350 ;
        RECT 135.955 201.960 136.835 202.130 ;
        RECT 137.670 201.440 137.930 203.090 ;
        RECT 154.660 202.450 155.540 202.620 ;
        RECT 154.240 202.230 154.410 202.400 ;
        RECT 155.790 202.230 155.960 202.400 ;
        RECT 154.660 202.010 155.540 202.180 ;
        RECT 158.005 202.460 158.885 202.630 ;
        RECT 157.540 202.240 157.710 202.410 ;
        RECT 159.180 202.240 159.350 202.410 ;
        RECT 158.005 202.020 158.885 202.190 ;
        RECT 159.720 201.500 159.980 203.150 ;
        RECT 132.610 200.290 133.490 200.460 ;
        RECT 132.190 200.070 132.360 200.240 ;
        RECT 133.740 200.070 133.910 200.240 ;
        RECT 132.610 199.850 133.490 200.020 ;
        RECT 135.955 200.300 136.835 200.470 ;
        RECT 135.490 200.080 135.660 200.250 ;
        RECT 137.130 200.080 137.300 200.250 ;
        RECT 135.955 199.860 136.835 200.030 ;
        RECT 137.670 199.340 137.930 200.990 ;
        RECT 154.660 200.350 155.540 200.520 ;
        RECT 154.240 200.130 154.410 200.300 ;
        RECT 155.790 200.130 155.960 200.300 ;
        RECT 154.660 199.910 155.540 200.080 ;
        RECT 158.005 200.360 158.885 200.530 ;
        RECT 157.540 200.140 157.710 200.310 ;
        RECT 159.180 200.140 159.350 200.310 ;
        RECT 158.005 199.920 158.885 200.090 ;
        RECT 159.720 199.400 159.980 201.050 ;
        RECT 132.610 198.200 133.490 198.370 ;
        RECT 132.190 197.980 132.360 198.150 ;
        RECT 133.740 197.980 133.910 198.150 ;
        RECT 132.610 197.760 133.490 197.930 ;
        RECT 135.955 198.210 136.835 198.380 ;
        RECT 135.490 197.990 135.660 198.160 ;
        RECT 137.130 197.990 137.300 198.160 ;
        RECT 135.955 197.770 136.835 197.940 ;
        RECT 137.670 197.250 137.930 198.900 ;
        RECT 154.660 198.250 155.540 198.420 ;
        RECT 154.240 198.030 154.410 198.200 ;
        RECT 155.790 198.030 155.960 198.200 ;
        RECT 154.660 197.810 155.540 197.980 ;
        RECT 158.005 198.260 158.885 198.430 ;
        RECT 157.540 198.040 157.710 198.210 ;
        RECT 159.180 198.040 159.350 198.210 ;
        RECT 158.005 197.820 158.885 197.990 ;
        RECT 159.720 197.300 159.980 198.950 ;
        RECT 132.610 196.100 133.490 196.270 ;
        RECT 132.190 195.880 132.360 196.050 ;
        RECT 133.740 195.880 133.910 196.050 ;
        RECT 132.610 195.660 133.490 195.830 ;
        RECT 135.955 196.110 136.835 196.280 ;
        RECT 135.490 195.890 135.660 196.060 ;
        RECT 137.130 195.890 137.300 196.060 ;
        RECT 135.955 195.670 136.835 195.840 ;
        RECT 137.670 195.150 137.930 196.800 ;
        RECT 154.660 196.150 155.540 196.320 ;
        RECT 154.240 195.930 154.410 196.100 ;
        RECT 155.790 195.930 155.960 196.100 ;
        RECT 154.660 195.710 155.540 195.880 ;
        RECT 158.005 196.160 158.885 196.330 ;
        RECT 157.540 195.940 157.710 196.110 ;
        RECT 159.180 195.940 159.350 196.110 ;
        RECT 158.005 195.720 158.885 195.890 ;
        RECT 159.720 195.200 159.980 196.850 ;
        RECT 132.610 194.000 133.490 194.170 ;
        RECT 132.190 193.780 132.360 193.950 ;
        RECT 133.740 193.780 133.910 193.950 ;
        RECT 132.610 193.560 133.490 193.730 ;
        RECT 135.955 194.010 136.835 194.180 ;
        RECT 135.490 193.790 135.660 193.960 ;
        RECT 137.130 193.790 137.300 193.960 ;
        RECT 135.955 193.570 136.835 193.740 ;
        RECT 137.670 193.050 137.930 194.700 ;
        RECT 154.660 194.050 155.540 194.220 ;
        RECT 154.240 193.830 154.410 194.000 ;
        RECT 155.790 193.830 155.960 194.000 ;
        RECT 154.660 193.610 155.540 193.780 ;
        RECT 158.005 194.060 158.885 194.230 ;
        RECT 157.540 193.840 157.710 194.010 ;
        RECT 159.180 193.840 159.350 194.010 ;
        RECT 158.005 193.620 158.885 193.790 ;
        RECT 159.720 193.100 159.980 194.750 ;
        RECT 132.610 191.900 133.490 192.070 ;
        RECT 132.190 191.680 132.360 191.850 ;
        RECT 133.740 191.680 133.910 191.850 ;
        RECT 132.610 191.460 133.490 191.630 ;
        RECT 135.955 191.910 136.835 192.080 ;
        RECT 135.490 191.690 135.660 191.860 ;
        RECT 137.130 191.690 137.300 191.860 ;
        RECT 135.955 191.470 136.835 191.640 ;
        RECT 137.670 190.950 137.930 192.600 ;
        RECT 154.660 191.950 155.540 192.120 ;
        RECT 154.240 191.730 154.410 191.900 ;
        RECT 155.790 191.730 155.960 191.900 ;
        RECT 154.660 191.510 155.540 191.680 ;
        RECT 158.005 191.960 158.885 192.130 ;
        RECT 157.540 191.740 157.710 191.910 ;
        RECT 159.180 191.740 159.350 191.910 ;
        RECT 158.005 191.520 158.885 191.690 ;
        RECT 159.720 191.000 159.980 192.650 ;
        RECT 132.610 189.800 133.490 189.970 ;
        RECT 132.190 189.580 132.360 189.750 ;
        RECT 133.740 189.580 133.910 189.750 ;
        RECT 132.610 189.360 133.490 189.530 ;
        RECT 135.955 189.810 136.835 189.980 ;
        RECT 135.490 189.590 135.660 189.760 ;
        RECT 137.130 189.590 137.300 189.760 ;
        RECT 135.955 189.370 136.835 189.540 ;
        RECT 137.670 188.850 137.930 190.500 ;
        RECT 154.660 189.850 155.540 190.020 ;
        RECT 154.240 189.630 154.410 189.800 ;
        RECT 155.790 189.630 155.960 189.800 ;
        RECT 154.660 189.410 155.540 189.580 ;
        RECT 158.005 189.860 158.885 190.030 ;
        RECT 157.540 189.640 157.710 189.810 ;
        RECT 159.180 189.640 159.350 189.810 ;
        RECT 158.005 189.420 158.885 189.590 ;
        RECT 159.720 188.900 159.980 190.550 ;
        RECT 132.610 187.700 133.490 187.870 ;
        RECT 132.190 187.480 132.360 187.650 ;
        RECT 133.740 187.480 133.910 187.650 ;
        RECT 132.610 187.260 133.490 187.430 ;
        RECT 135.955 187.710 136.835 187.880 ;
        RECT 135.490 187.490 135.660 187.660 ;
        RECT 137.130 187.490 137.300 187.660 ;
        RECT 135.955 187.270 136.835 187.440 ;
        RECT 137.670 186.750 137.930 188.400 ;
        RECT 154.660 187.750 155.540 187.920 ;
        RECT 154.240 187.530 154.410 187.700 ;
        RECT 155.790 187.530 155.960 187.700 ;
        RECT 154.660 187.310 155.540 187.480 ;
        RECT 158.005 187.760 158.885 187.930 ;
        RECT 157.540 187.540 157.710 187.710 ;
        RECT 159.180 187.540 159.350 187.710 ;
        RECT 158.005 187.320 158.885 187.490 ;
        RECT 159.720 186.800 159.980 188.450 ;
        RECT 132.610 185.600 133.490 185.770 ;
        RECT 132.190 185.380 132.360 185.550 ;
        RECT 133.740 185.380 133.910 185.550 ;
        RECT 132.610 185.160 133.490 185.330 ;
        RECT 135.955 185.610 136.835 185.780 ;
        RECT 135.490 185.390 135.660 185.560 ;
        RECT 137.130 185.390 137.300 185.560 ;
        RECT 135.955 185.170 136.835 185.340 ;
        RECT 137.670 184.650 137.930 186.300 ;
        RECT 154.660 185.650 155.540 185.820 ;
        RECT 154.240 185.430 154.410 185.600 ;
        RECT 155.790 185.430 155.960 185.600 ;
        RECT 154.660 185.210 155.540 185.380 ;
        RECT 158.005 185.660 158.885 185.830 ;
        RECT 157.540 185.440 157.710 185.610 ;
        RECT 159.180 185.440 159.350 185.610 ;
        RECT 158.005 185.220 158.885 185.390 ;
        RECT 159.720 184.700 159.980 186.350 ;
        RECT 132.610 183.500 133.490 183.670 ;
        RECT 132.190 183.280 132.360 183.450 ;
        RECT 133.740 183.280 133.910 183.450 ;
        RECT 132.610 183.060 133.490 183.230 ;
        RECT 135.955 183.510 136.835 183.680 ;
        RECT 135.490 183.290 135.660 183.460 ;
        RECT 137.130 183.290 137.300 183.460 ;
        RECT 135.955 183.070 136.835 183.240 ;
        RECT 137.670 182.550 137.930 184.200 ;
        RECT 154.660 183.550 155.540 183.720 ;
        RECT 154.240 183.330 154.410 183.500 ;
        RECT 155.790 183.330 155.960 183.500 ;
        RECT 154.660 183.110 155.540 183.280 ;
        RECT 158.005 183.560 158.885 183.730 ;
        RECT 157.540 183.340 157.710 183.510 ;
        RECT 159.180 183.340 159.350 183.510 ;
        RECT 158.005 183.120 158.885 183.290 ;
        RECT 159.720 182.600 159.980 184.250 ;
        RECT 132.610 181.400 133.490 181.570 ;
        RECT 132.190 181.180 132.360 181.350 ;
        RECT 133.740 181.180 133.910 181.350 ;
        RECT 132.610 180.960 133.490 181.130 ;
        RECT 135.955 181.410 136.835 181.580 ;
        RECT 135.490 181.190 135.660 181.360 ;
        RECT 137.130 181.190 137.300 181.360 ;
        RECT 135.955 180.970 136.835 181.140 ;
        RECT 137.670 180.450 137.930 182.100 ;
        RECT 154.660 181.450 155.540 181.620 ;
        RECT 154.240 181.230 154.410 181.400 ;
        RECT 155.790 181.230 155.960 181.400 ;
        RECT 154.660 181.010 155.540 181.180 ;
        RECT 158.005 181.460 158.885 181.630 ;
        RECT 157.540 181.240 157.710 181.410 ;
        RECT 159.180 181.240 159.350 181.410 ;
        RECT 158.005 181.020 158.885 181.190 ;
        RECT 159.720 180.500 159.980 182.150 ;
        RECT 132.610 179.310 133.490 179.480 ;
        RECT 132.190 179.090 132.360 179.260 ;
        RECT 133.740 179.090 133.910 179.260 ;
        RECT 132.610 178.870 133.490 179.040 ;
        RECT 135.955 179.320 136.835 179.490 ;
        RECT 135.490 179.100 135.660 179.270 ;
        RECT 137.130 179.100 137.300 179.270 ;
        RECT 135.955 178.880 136.835 179.050 ;
        RECT 137.670 178.360 137.930 180.010 ;
        RECT 154.660 179.350 155.540 179.520 ;
        RECT 154.240 179.130 154.410 179.300 ;
        RECT 155.790 179.130 155.960 179.300 ;
        RECT 154.660 178.910 155.540 179.080 ;
        RECT 158.005 179.360 158.885 179.530 ;
        RECT 157.540 179.140 157.710 179.310 ;
        RECT 159.180 179.140 159.350 179.310 ;
        RECT 158.005 178.920 158.885 179.090 ;
        RECT 159.720 178.400 159.980 180.050 ;
        RECT 132.610 177.220 133.490 177.390 ;
        RECT 132.190 177.000 132.360 177.170 ;
        RECT 133.740 177.000 133.910 177.170 ;
        RECT 132.610 176.780 133.490 176.950 ;
        RECT 135.955 177.230 136.835 177.400 ;
        RECT 135.490 177.010 135.660 177.180 ;
        RECT 137.130 177.010 137.300 177.180 ;
        RECT 135.955 176.790 136.835 176.960 ;
        RECT 137.670 176.270 137.930 177.920 ;
        RECT 154.660 177.250 155.540 177.420 ;
        RECT 154.240 177.030 154.410 177.200 ;
        RECT 155.790 177.030 155.960 177.200 ;
        RECT 154.660 176.810 155.540 176.980 ;
        RECT 158.005 177.260 158.885 177.430 ;
        RECT 157.540 177.040 157.710 177.210 ;
        RECT 159.180 177.040 159.350 177.210 ;
        RECT 158.005 176.820 158.885 176.990 ;
        RECT 159.720 176.300 159.980 177.950 ;
        RECT 132.610 175.120 133.490 175.290 ;
        RECT 132.190 174.900 132.360 175.070 ;
        RECT 133.740 174.900 133.910 175.070 ;
        RECT 132.610 174.680 133.490 174.850 ;
        RECT 135.955 175.130 136.835 175.300 ;
        RECT 135.490 174.910 135.660 175.080 ;
        RECT 137.130 174.910 137.300 175.080 ;
        RECT 135.955 174.690 136.835 174.860 ;
        RECT 137.670 174.170 137.930 175.820 ;
        RECT 154.660 175.150 155.540 175.320 ;
        RECT 154.240 174.930 154.410 175.100 ;
        RECT 155.790 174.930 155.960 175.100 ;
        RECT 154.660 174.710 155.540 174.880 ;
        RECT 158.005 175.160 158.885 175.330 ;
        RECT 157.540 174.940 157.710 175.110 ;
        RECT 159.180 174.940 159.350 175.110 ;
        RECT 158.005 174.720 158.885 174.890 ;
        RECT 159.720 174.200 159.980 175.850 ;
        RECT 132.610 173.030 133.490 173.200 ;
        RECT 132.190 172.810 132.360 172.980 ;
        RECT 133.740 172.810 133.910 172.980 ;
        RECT 132.610 172.590 133.490 172.760 ;
        RECT 135.955 173.040 136.835 173.210 ;
        RECT 135.490 172.820 135.660 172.990 ;
        RECT 137.130 172.820 137.300 172.990 ;
        RECT 135.955 172.600 136.835 172.770 ;
        RECT 137.670 172.080 137.930 173.730 ;
        RECT 154.660 173.050 155.540 173.220 ;
        RECT 154.240 172.830 154.410 173.000 ;
        RECT 155.790 172.830 155.960 173.000 ;
        RECT 154.660 172.610 155.540 172.780 ;
        RECT 158.005 173.060 158.885 173.230 ;
        RECT 157.540 172.840 157.710 173.010 ;
        RECT 159.180 172.840 159.350 173.010 ;
        RECT 158.005 172.620 158.885 172.790 ;
        RECT 159.720 172.100 159.980 173.750 ;
        RECT 132.610 170.940 133.490 171.110 ;
        RECT 132.190 170.720 132.360 170.890 ;
        RECT 133.740 170.720 133.910 170.890 ;
        RECT 132.610 170.500 133.490 170.670 ;
        RECT 135.955 170.950 136.835 171.120 ;
        RECT 135.490 170.730 135.660 170.900 ;
        RECT 137.130 170.730 137.300 170.900 ;
        RECT 135.955 170.510 136.835 170.680 ;
        RECT 137.670 169.990 137.930 171.640 ;
        RECT 154.660 170.950 155.540 171.120 ;
        RECT 154.240 170.730 154.410 170.900 ;
        RECT 155.790 170.730 155.960 170.900 ;
        RECT 154.660 170.510 155.540 170.680 ;
        RECT 158.005 170.960 158.885 171.130 ;
        RECT 157.540 170.740 157.710 170.910 ;
        RECT 159.180 170.740 159.350 170.910 ;
        RECT 158.005 170.520 158.885 170.690 ;
        RECT 159.720 170.000 159.980 171.650 ;
        RECT 132.610 168.840 133.490 169.010 ;
        RECT 132.190 168.620 132.360 168.790 ;
        RECT 133.740 168.620 133.910 168.790 ;
        RECT 132.610 168.400 133.490 168.570 ;
        RECT 135.955 168.850 136.835 169.020 ;
        RECT 135.490 168.630 135.660 168.800 ;
        RECT 137.130 168.630 137.300 168.800 ;
        RECT 135.955 168.410 136.835 168.580 ;
        RECT 137.670 167.890 137.930 169.540 ;
        RECT 154.660 168.850 155.540 169.020 ;
        RECT 154.240 168.630 154.410 168.800 ;
        RECT 155.790 168.630 155.960 168.800 ;
        RECT 154.660 168.410 155.540 168.580 ;
        RECT 158.005 168.860 158.885 169.030 ;
        RECT 157.540 168.640 157.710 168.810 ;
        RECT 159.180 168.640 159.350 168.810 ;
        RECT 158.005 168.420 158.885 168.590 ;
        RECT 159.720 167.900 159.980 169.550 ;
        RECT 132.610 166.740 133.490 166.910 ;
        RECT 132.190 166.520 132.360 166.690 ;
        RECT 133.740 166.520 133.910 166.690 ;
        RECT 132.610 166.300 133.490 166.470 ;
        RECT 135.955 166.750 136.835 166.920 ;
        RECT 135.490 166.530 135.660 166.700 ;
        RECT 137.130 166.530 137.300 166.700 ;
        RECT 135.955 166.310 136.835 166.480 ;
        RECT 137.670 165.790 137.930 167.440 ;
        RECT 154.660 166.750 155.540 166.920 ;
        RECT 154.240 166.530 154.410 166.700 ;
        RECT 155.790 166.530 155.960 166.700 ;
        RECT 154.660 166.310 155.540 166.480 ;
        RECT 158.005 166.760 158.885 166.930 ;
        RECT 157.540 166.540 157.710 166.710 ;
        RECT 159.180 166.540 159.350 166.710 ;
        RECT 158.005 166.320 158.885 166.490 ;
        RECT 159.720 165.800 159.980 167.450 ;
        RECT 132.610 164.640 133.490 164.810 ;
        RECT 132.190 164.420 132.360 164.590 ;
        RECT 133.740 164.420 133.910 164.590 ;
        RECT 132.610 164.200 133.490 164.370 ;
        RECT 135.955 164.650 136.835 164.820 ;
        RECT 135.490 164.430 135.660 164.600 ;
        RECT 137.130 164.430 137.300 164.600 ;
        RECT 135.955 164.210 136.835 164.380 ;
        RECT 137.670 163.690 137.930 165.340 ;
        RECT 154.660 164.650 155.540 164.820 ;
        RECT 154.240 164.430 154.410 164.600 ;
        RECT 155.790 164.430 155.960 164.600 ;
        RECT 154.660 164.210 155.540 164.380 ;
        RECT 158.005 164.660 158.885 164.830 ;
        RECT 157.540 164.440 157.710 164.610 ;
        RECT 159.180 164.440 159.350 164.610 ;
        RECT 158.005 164.220 158.885 164.390 ;
        RECT 159.720 163.700 159.980 165.350 ;
        RECT 132.610 162.540 133.490 162.710 ;
        RECT 132.190 162.320 132.360 162.490 ;
        RECT 133.740 162.320 133.910 162.490 ;
        RECT 132.610 162.100 133.490 162.270 ;
        RECT 135.955 162.550 136.835 162.720 ;
        RECT 135.490 162.330 135.660 162.500 ;
        RECT 137.130 162.330 137.300 162.500 ;
        RECT 135.955 162.110 136.835 162.280 ;
        RECT 137.670 161.590 137.930 163.240 ;
        RECT 154.660 162.550 155.540 162.720 ;
        RECT 154.240 162.330 154.410 162.500 ;
        RECT 155.790 162.330 155.960 162.500 ;
        RECT 154.660 162.110 155.540 162.280 ;
        RECT 158.005 162.560 158.885 162.730 ;
        RECT 157.540 162.340 157.710 162.510 ;
        RECT 159.180 162.340 159.350 162.510 ;
        RECT 158.005 162.120 158.885 162.290 ;
        RECT 159.720 161.600 159.980 163.250 ;
        RECT 132.610 160.440 133.490 160.610 ;
        RECT 132.190 160.220 132.360 160.390 ;
        RECT 133.740 160.220 133.910 160.390 ;
        RECT 132.610 160.000 133.490 160.170 ;
        RECT 135.955 160.450 136.835 160.620 ;
        RECT 135.490 160.230 135.660 160.400 ;
        RECT 137.130 160.230 137.300 160.400 ;
        RECT 135.955 160.010 136.835 160.180 ;
        RECT 137.670 159.490 137.930 161.140 ;
        RECT 154.660 160.450 155.540 160.620 ;
        RECT 154.240 160.230 154.410 160.400 ;
        RECT 155.790 160.230 155.960 160.400 ;
        RECT 154.660 160.010 155.540 160.180 ;
        RECT 158.005 160.460 158.885 160.630 ;
        RECT 157.540 160.240 157.710 160.410 ;
        RECT 159.180 160.240 159.350 160.410 ;
        RECT 158.005 160.020 158.885 160.190 ;
        RECT 159.720 159.500 159.980 161.150 ;
        RECT 132.610 158.340 133.490 158.510 ;
        RECT 132.190 158.120 132.360 158.290 ;
        RECT 133.740 158.120 133.910 158.290 ;
        RECT 132.610 157.900 133.490 158.070 ;
        RECT 135.955 158.350 136.835 158.520 ;
        RECT 135.490 158.130 135.660 158.300 ;
        RECT 137.130 158.130 137.300 158.300 ;
        RECT 135.955 157.910 136.835 158.080 ;
        RECT 137.670 157.390 137.930 159.040 ;
        RECT 154.660 158.350 155.540 158.520 ;
        RECT 154.240 158.130 154.410 158.300 ;
        RECT 155.790 158.130 155.960 158.300 ;
        RECT 154.660 157.910 155.540 158.080 ;
        RECT 158.005 158.360 158.885 158.530 ;
        RECT 157.540 158.140 157.710 158.310 ;
        RECT 159.180 158.140 159.350 158.310 ;
        RECT 158.005 157.920 158.885 158.090 ;
        RECT 159.720 157.400 159.980 159.050 ;
        RECT 132.610 156.240 133.490 156.410 ;
        RECT 132.190 156.020 132.360 156.190 ;
        RECT 133.740 156.020 133.910 156.190 ;
        RECT 132.610 155.800 133.490 155.970 ;
        RECT 135.955 156.250 136.835 156.420 ;
        RECT 135.490 156.030 135.660 156.200 ;
        RECT 137.130 156.030 137.300 156.200 ;
        RECT 135.955 155.810 136.835 155.980 ;
        RECT 137.670 155.290 137.930 156.940 ;
        RECT 154.660 156.250 155.540 156.420 ;
        RECT 154.240 156.030 154.410 156.200 ;
        RECT 155.790 156.030 155.960 156.200 ;
        RECT 154.660 155.810 155.540 155.980 ;
        RECT 158.005 156.260 158.885 156.430 ;
        RECT 157.540 156.040 157.710 156.210 ;
        RECT 159.180 156.040 159.350 156.210 ;
        RECT 158.005 155.820 158.885 155.990 ;
        RECT 159.720 155.300 159.980 156.950 ;
        RECT 132.610 154.140 133.490 154.310 ;
        RECT 132.190 153.920 132.360 154.090 ;
        RECT 133.740 153.920 133.910 154.090 ;
        RECT 132.610 153.700 133.490 153.870 ;
        RECT 135.955 154.150 136.835 154.320 ;
        RECT 135.490 153.930 135.660 154.100 ;
        RECT 137.130 153.930 137.300 154.100 ;
        RECT 135.955 153.710 136.835 153.880 ;
        RECT 137.670 153.190 137.930 154.840 ;
        RECT 154.660 154.150 155.540 154.320 ;
        RECT 154.240 153.930 154.410 154.100 ;
        RECT 155.790 153.930 155.960 154.100 ;
        RECT 154.660 153.710 155.540 153.880 ;
        RECT 158.005 154.160 158.885 154.330 ;
        RECT 157.540 153.940 157.710 154.110 ;
        RECT 159.180 153.940 159.350 154.110 ;
        RECT 158.005 153.720 158.885 153.890 ;
        RECT 159.720 153.200 159.980 154.850 ;
        RECT 132.610 152.040 133.490 152.210 ;
        RECT 132.190 151.820 132.360 151.990 ;
        RECT 133.740 151.820 133.910 151.990 ;
        RECT 132.610 151.600 133.490 151.770 ;
        RECT 135.955 152.050 136.835 152.220 ;
        RECT 135.490 151.830 135.660 152.000 ;
        RECT 137.130 151.830 137.300 152.000 ;
        RECT 135.955 151.610 136.835 151.780 ;
        RECT 137.670 151.090 137.930 152.740 ;
        RECT 154.660 152.050 155.540 152.220 ;
        RECT 154.240 151.830 154.410 152.000 ;
        RECT 155.790 151.830 155.960 152.000 ;
        RECT 154.660 151.610 155.540 151.780 ;
        RECT 158.005 152.060 158.885 152.230 ;
        RECT 157.540 151.840 157.710 152.010 ;
        RECT 159.180 151.840 159.350 152.010 ;
        RECT 158.005 151.620 158.885 151.790 ;
        RECT 159.720 151.100 159.980 152.750 ;
        RECT 132.610 149.940 133.490 150.110 ;
        RECT 132.190 149.720 132.360 149.890 ;
        RECT 133.740 149.720 133.910 149.890 ;
        RECT 132.610 149.500 133.490 149.670 ;
        RECT 135.955 149.950 136.835 150.120 ;
        RECT 135.490 149.730 135.660 149.900 ;
        RECT 137.130 149.730 137.300 149.900 ;
        RECT 135.955 149.510 136.835 149.680 ;
        RECT 137.670 148.990 137.930 150.640 ;
        RECT 154.660 149.950 155.540 150.120 ;
        RECT 154.240 149.730 154.410 149.900 ;
        RECT 155.790 149.730 155.960 149.900 ;
        RECT 154.660 149.510 155.540 149.680 ;
        RECT 158.005 149.960 158.885 150.130 ;
        RECT 157.540 149.740 157.710 149.910 ;
        RECT 159.180 149.740 159.350 149.910 ;
        RECT 158.005 149.520 158.885 149.690 ;
        RECT 159.720 149.000 159.980 150.650 ;
        RECT 132.610 147.840 133.490 148.010 ;
        RECT 132.190 147.620 132.360 147.790 ;
        RECT 133.740 147.620 133.910 147.790 ;
        RECT 132.610 147.400 133.490 147.570 ;
        RECT 135.955 147.850 136.835 148.020 ;
        RECT 135.490 147.630 135.660 147.800 ;
        RECT 137.130 147.630 137.300 147.800 ;
        RECT 135.955 147.410 136.835 147.580 ;
        RECT 137.670 146.890 137.930 148.540 ;
        RECT 154.660 147.850 155.540 148.020 ;
        RECT 154.240 147.630 154.410 147.800 ;
        RECT 155.790 147.630 155.960 147.800 ;
        RECT 154.660 147.410 155.540 147.580 ;
        RECT 158.005 147.860 158.885 148.030 ;
        RECT 157.540 147.640 157.710 147.810 ;
        RECT 159.180 147.640 159.350 147.810 ;
        RECT 158.005 147.420 158.885 147.590 ;
        RECT 159.720 146.900 159.980 148.550 ;
        RECT 132.610 145.740 133.490 145.910 ;
        RECT 132.190 145.520 132.360 145.690 ;
        RECT 133.740 145.520 133.910 145.690 ;
        RECT 132.610 145.300 133.490 145.470 ;
        RECT 135.955 145.750 136.835 145.920 ;
        RECT 135.490 145.530 135.660 145.700 ;
        RECT 137.130 145.530 137.300 145.700 ;
        RECT 135.955 145.310 136.835 145.480 ;
        RECT 137.670 144.790 137.930 146.440 ;
        RECT 154.660 145.750 155.540 145.920 ;
        RECT 154.240 145.530 154.410 145.700 ;
        RECT 155.790 145.530 155.960 145.700 ;
        RECT 154.660 145.310 155.540 145.480 ;
        RECT 158.005 145.760 158.885 145.930 ;
        RECT 157.540 145.540 157.710 145.710 ;
        RECT 159.180 145.540 159.350 145.710 ;
        RECT 158.005 145.320 158.885 145.490 ;
        RECT 159.720 144.800 159.980 146.450 ;
        RECT 132.610 143.640 133.490 143.810 ;
        RECT 132.190 143.420 132.360 143.590 ;
        RECT 133.740 143.420 133.910 143.590 ;
        RECT 132.610 143.200 133.490 143.370 ;
        RECT 135.955 143.650 136.835 143.820 ;
        RECT 135.490 143.430 135.660 143.600 ;
        RECT 137.130 143.430 137.300 143.600 ;
        RECT 135.955 143.210 136.835 143.380 ;
        RECT 137.670 142.690 137.930 144.340 ;
        RECT 154.660 143.650 155.540 143.820 ;
        RECT 154.240 143.430 154.410 143.600 ;
        RECT 155.790 143.430 155.960 143.600 ;
        RECT 154.660 143.210 155.540 143.380 ;
        RECT 158.005 143.660 158.885 143.830 ;
        RECT 157.540 143.440 157.710 143.610 ;
        RECT 159.180 143.440 159.350 143.610 ;
        RECT 158.005 143.220 158.885 143.390 ;
        RECT 159.720 142.700 159.980 144.350 ;
        RECT 132.610 141.540 133.490 141.710 ;
        RECT 132.190 141.320 132.360 141.490 ;
        RECT 133.740 141.320 133.910 141.490 ;
        RECT 132.610 141.100 133.490 141.270 ;
        RECT 135.955 141.550 136.835 141.720 ;
        RECT 135.490 141.330 135.660 141.500 ;
        RECT 137.130 141.330 137.300 141.500 ;
        RECT 135.955 141.110 136.835 141.280 ;
        RECT 137.670 140.590 137.930 142.240 ;
        RECT 154.660 141.550 155.540 141.720 ;
        RECT 154.240 141.330 154.410 141.500 ;
        RECT 155.790 141.330 155.960 141.500 ;
        RECT 154.660 141.110 155.540 141.280 ;
        RECT 158.005 141.560 158.885 141.730 ;
        RECT 157.540 141.340 157.710 141.510 ;
        RECT 159.180 141.340 159.350 141.510 ;
        RECT 158.005 141.120 158.885 141.290 ;
        RECT 159.720 140.600 159.980 142.250 ;
        RECT 132.610 139.440 133.490 139.610 ;
        RECT 132.190 139.220 132.360 139.390 ;
        RECT 133.740 139.220 133.910 139.390 ;
        RECT 132.610 139.000 133.490 139.170 ;
        RECT 135.955 139.450 136.835 139.620 ;
        RECT 135.490 139.230 135.660 139.400 ;
        RECT 137.130 139.230 137.300 139.400 ;
        RECT 135.955 139.010 136.835 139.180 ;
        RECT 137.670 138.490 137.930 140.140 ;
        RECT 154.660 139.450 155.540 139.620 ;
        RECT 154.240 139.230 154.410 139.400 ;
        RECT 155.790 139.230 155.960 139.400 ;
        RECT 154.660 139.010 155.540 139.180 ;
        RECT 158.005 139.460 158.885 139.630 ;
        RECT 157.540 139.240 157.710 139.410 ;
        RECT 159.180 139.240 159.350 139.410 ;
        RECT 158.005 139.020 158.885 139.190 ;
        RECT 159.720 138.500 159.980 140.150 ;
        RECT 132.610 137.340 133.490 137.510 ;
        RECT 132.190 137.120 132.360 137.290 ;
        RECT 133.740 137.120 133.910 137.290 ;
        RECT 132.610 136.900 133.490 137.070 ;
        RECT 135.955 137.350 136.835 137.520 ;
        RECT 135.490 137.130 135.660 137.300 ;
        RECT 137.130 137.130 137.300 137.300 ;
        RECT 135.955 136.910 136.835 137.080 ;
        RECT 137.670 136.390 137.930 138.040 ;
        RECT 154.660 137.350 155.540 137.520 ;
        RECT 154.240 137.130 154.410 137.300 ;
        RECT 155.790 137.130 155.960 137.300 ;
        RECT 154.660 136.910 155.540 137.080 ;
        RECT 158.005 137.360 158.885 137.530 ;
        RECT 157.540 137.140 157.710 137.310 ;
        RECT 159.180 137.140 159.350 137.310 ;
        RECT 158.005 136.920 158.885 137.090 ;
        RECT 159.720 136.400 159.980 138.050 ;
        RECT 132.610 135.240 133.490 135.410 ;
        RECT 132.190 135.020 132.360 135.190 ;
        RECT 133.740 135.020 133.910 135.190 ;
        RECT 132.610 134.800 133.490 134.970 ;
        RECT 135.955 135.250 136.835 135.420 ;
        RECT 135.490 135.030 135.660 135.200 ;
        RECT 137.130 135.030 137.300 135.200 ;
        RECT 135.955 134.810 136.835 134.980 ;
        RECT 137.670 134.290 137.930 135.940 ;
        RECT 154.660 135.250 155.540 135.420 ;
        RECT 154.240 135.030 154.410 135.200 ;
        RECT 155.790 135.030 155.960 135.200 ;
        RECT 154.660 134.810 155.540 134.980 ;
        RECT 158.005 135.260 158.885 135.430 ;
        RECT 157.540 135.040 157.710 135.210 ;
        RECT 159.180 135.040 159.350 135.210 ;
        RECT 158.005 134.820 158.885 134.990 ;
        RECT 159.720 134.300 159.980 135.950 ;
        RECT 132.610 133.140 133.490 133.310 ;
        RECT 132.190 132.920 132.360 133.090 ;
        RECT 133.740 132.920 133.910 133.090 ;
        RECT 132.610 132.700 133.490 132.870 ;
        RECT 135.955 133.150 136.835 133.320 ;
        RECT 135.490 132.930 135.660 133.100 ;
        RECT 137.130 132.930 137.300 133.100 ;
        RECT 135.955 132.710 136.835 132.880 ;
        RECT 137.670 132.190 137.930 133.840 ;
        RECT 154.660 133.150 155.540 133.320 ;
        RECT 154.240 132.930 154.410 133.100 ;
        RECT 155.790 132.930 155.960 133.100 ;
        RECT 154.660 132.710 155.540 132.880 ;
        RECT 158.005 133.160 158.885 133.330 ;
        RECT 157.540 132.940 157.710 133.110 ;
        RECT 159.180 132.940 159.350 133.110 ;
        RECT 158.005 132.720 158.885 132.890 ;
        RECT 159.720 132.200 159.980 133.850 ;
        RECT 132.610 131.040 133.490 131.210 ;
        RECT 132.190 130.820 132.360 130.990 ;
        RECT 133.740 130.820 133.910 130.990 ;
        RECT 132.610 130.600 133.490 130.770 ;
        RECT 135.955 131.050 136.835 131.220 ;
        RECT 135.490 130.830 135.660 131.000 ;
        RECT 137.130 130.830 137.300 131.000 ;
        RECT 135.955 130.610 136.835 130.780 ;
        RECT 137.670 130.090 137.930 131.740 ;
        RECT 154.660 131.050 155.540 131.220 ;
        RECT 154.240 130.830 154.410 131.000 ;
        RECT 155.790 130.830 155.960 131.000 ;
        RECT 154.660 130.610 155.540 130.780 ;
        RECT 158.005 131.060 158.885 131.230 ;
        RECT 157.540 130.840 157.710 131.010 ;
        RECT 159.180 130.840 159.350 131.010 ;
        RECT 158.005 130.620 158.885 130.790 ;
        RECT 159.720 130.100 159.980 131.750 ;
        RECT 132.610 128.940 133.490 129.110 ;
        RECT 132.190 128.720 132.360 128.890 ;
        RECT 133.740 128.720 133.910 128.890 ;
        RECT 132.610 128.500 133.490 128.670 ;
        RECT 135.955 128.950 136.835 129.120 ;
        RECT 135.490 128.730 135.660 128.900 ;
        RECT 137.130 128.730 137.300 128.900 ;
        RECT 135.955 128.510 136.835 128.680 ;
        RECT 137.670 127.990 137.930 129.640 ;
        RECT 154.660 128.950 155.540 129.120 ;
        RECT 154.240 128.730 154.410 128.900 ;
        RECT 155.790 128.730 155.960 128.900 ;
        RECT 154.660 128.510 155.540 128.680 ;
        RECT 158.005 128.960 158.885 129.130 ;
        RECT 157.540 128.740 157.710 128.910 ;
        RECT 159.180 128.740 159.350 128.910 ;
        RECT 158.005 128.520 158.885 128.690 ;
        RECT 159.720 128.000 159.980 129.650 ;
        RECT 132.610 126.840 133.490 127.010 ;
        RECT 132.190 126.620 132.360 126.790 ;
        RECT 133.740 126.620 133.910 126.790 ;
        RECT 132.610 126.400 133.490 126.570 ;
        RECT 135.955 126.850 136.835 127.020 ;
        RECT 135.490 126.630 135.660 126.800 ;
        RECT 137.130 126.630 137.300 126.800 ;
        RECT 135.955 126.410 136.835 126.580 ;
        RECT 137.670 125.890 137.930 127.540 ;
        RECT 154.660 126.850 155.540 127.020 ;
        RECT 154.240 126.630 154.410 126.800 ;
        RECT 155.790 126.630 155.960 126.800 ;
        RECT 154.660 126.410 155.540 126.580 ;
        RECT 158.005 126.860 158.885 127.030 ;
        RECT 157.540 126.640 157.710 126.810 ;
        RECT 159.180 126.640 159.350 126.810 ;
        RECT 158.005 126.420 158.885 126.590 ;
        RECT 159.720 125.900 159.980 127.550 ;
        RECT 132.610 124.740 133.490 124.910 ;
        RECT 132.190 124.520 132.360 124.690 ;
        RECT 133.740 124.520 133.910 124.690 ;
        RECT 132.610 124.300 133.490 124.470 ;
        RECT 135.955 124.750 136.835 124.920 ;
        RECT 135.490 124.530 135.660 124.700 ;
        RECT 137.130 124.530 137.300 124.700 ;
        RECT 135.955 124.310 136.835 124.480 ;
        RECT 137.670 123.790 137.930 125.440 ;
        RECT 154.660 124.750 155.540 124.920 ;
        RECT 154.240 124.530 154.410 124.700 ;
        RECT 155.790 124.530 155.960 124.700 ;
        RECT 154.660 124.310 155.540 124.480 ;
        RECT 158.005 124.760 158.885 124.930 ;
        RECT 157.540 124.540 157.710 124.710 ;
        RECT 159.180 124.540 159.350 124.710 ;
        RECT 158.005 124.320 158.885 124.490 ;
        RECT 159.720 123.800 159.980 125.450 ;
        RECT 132.610 122.640 133.490 122.810 ;
        RECT 132.190 122.420 132.360 122.590 ;
        RECT 133.740 122.420 133.910 122.590 ;
        RECT 132.610 122.200 133.490 122.370 ;
        RECT 135.955 122.650 136.835 122.820 ;
        RECT 135.490 122.430 135.660 122.600 ;
        RECT 137.130 122.430 137.300 122.600 ;
        RECT 135.955 122.210 136.835 122.380 ;
        RECT 137.670 121.690 137.930 123.340 ;
        RECT 154.660 122.650 155.540 122.820 ;
        RECT 154.240 122.430 154.410 122.600 ;
        RECT 155.790 122.430 155.960 122.600 ;
        RECT 154.660 122.210 155.540 122.380 ;
        RECT 158.005 122.660 158.885 122.830 ;
        RECT 157.540 122.440 157.710 122.610 ;
        RECT 159.180 122.440 159.350 122.610 ;
        RECT 158.005 122.220 158.885 122.390 ;
        RECT 159.720 121.700 159.980 123.350 ;
        RECT 132.610 120.540 133.490 120.710 ;
        RECT 132.190 120.320 132.360 120.490 ;
        RECT 133.740 120.320 133.910 120.490 ;
        RECT 132.610 120.100 133.490 120.270 ;
        RECT 135.955 120.550 136.835 120.720 ;
        RECT 135.490 120.330 135.660 120.500 ;
        RECT 137.130 120.330 137.300 120.500 ;
        RECT 135.955 120.110 136.835 120.280 ;
        RECT 137.670 119.590 137.930 121.240 ;
        RECT 154.660 120.550 155.540 120.720 ;
        RECT 154.240 120.330 154.410 120.500 ;
        RECT 155.790 120.330 155.960 120.500 ;
        RECT 154.660 120.110 155.540 120.280 ;
        RECT 158.005 120.560 158.885 120.730 ;
        RECT 157.540 120.340 157.710 120.510 ;
        RECT 159.180 120.340 159.350 120.510 ;
        RECT 158.005 120.120 158.885 120.290 ;
        RECT 159.720 119.600 159.980 121.250 ;
        RECT 132.610 118.440 133.490 118.610 ;
        RECT 132.190 118.220 132.360 118.390 ;
        RECT 133.740 118.220 133.910 118.390 ;
        RECT 132.610 118.000 133.490 118.170 ;
        RECT 135.955 118.450 136.835 118.620 ;
        RECT 135.490 118.230 135.660 118.400 ;
        RECT 137.130 118.230 137.300 118.400 ;
        RECT 135.955 118.010 136.835 118.180 ;
        RECT 137.670 117.490 137.930 119.140 ;
        RECT 154.660 118.450 155.540 118.620 ;
        RECT 154.240 118.230 154.410 118.400 ;
        RECT 155.790 118.230 155.960 118.400 ;
        RECT 154.660 118.010 155.540 118.180 ;
        RECT 158.005 118.460 158.885 118.630 ;
        RECT 157.540 118.240 157.710 118.410 ;
        RECT 159.180 118.240 159.350 118.410 ;
        RECT 158.005 118.020 158.885 118.190 ;
        RECT 159.720 117.500 159.980 119.150 ;
        RECT 132.610 116.340 133.490 116.510 ;
        RECT 132.190 116.120 132.360 116.290 ;
        RECT 133.740 116.120 133.910 116.290 ;
        RECT 132.610 115.900 133.490 116.070 ;
        RECT 135.955 116.350 136.835 116.520 ;
        RECT 135.490 116.130 135.660 116.300 ;
        RECT 137.130 116.130 137.300 116.300 ;
        RECT 135.955 115.910 136.835 116.080 ;
        RECT 137.670 115.390 137.930 117.040 ;
        RECT 154.660 116.350 155.540 116.520 ;
        RECT 154.240 116.130 154.410 116.300 ;
        RECT 155.790 116.130 155.960 116.300 ;
        RECT 154.660 115.910 155.540 116.080 ;
        RECT 158.005 116.360 158.885 116.530 ;
        RECT 157.540 116.140 157.710 116.310 ;
        RECT 159.180 116.140 159.350 116.310 ;
        RECT 158.005 115.920 158.885 116.090 ;
        RECT 159.720 115.400 159.980 117.050 ;
        RECT 132.610 114.240 133.490 114.410 ;
        RECT 132.190 114.020 132.360 114.190 ;
        RECT 133.740 114.020 133.910 114.190 ;
        RECT 132.610 113.800 133.490 113.970 ;
        RECT 135.955 114.250 136.835 114.420 ;
        RECT 135.490 114.030 135.660 114.200 ;
        RECT 137.130 114.030 137.300 114.200 ;
        RECT 135.955 113.810 136.835 113.980 ;
        RECT 137.670 113.290 137.930 114.940 ;
        RECT 154.660 114.250 155.540 114.420 ;
        RECT 154.240 114.030 154.410 114.200 ;
        RECT 155.790 114.030 155.960 114.200 ;
        RECT 154.660 113.810 155.540 113.980 ;
        RECT 158.005 114.260 158.885 114.430 ;
        RECT 157.540 114.040 157.710 114.210 ;
        RECT 159.180 114.040 159.350 114.210 ;
        RECT 158.005 113.820 158.885 113.990 ;
        RECT 159.720 113.300 159.980 114.950 ;
        RECT 132.610 112.140 133.490 112.310 ;
        RECT 132.190 111.920 132.360 112.090 ;
        RECT 133.740 111.920 133.910 112.090 ;
        RECT 132.610 111.700 133.490 111.870 ;
        RECT 135.955 112.150 136.835 112.320 ;
        RECT 135.490 111.930 135.660 112.100 ;
        RECT 137.130 111.930 137.300 112.100 ;
        RECT 135.955 111.710 136.835 111.880 ;
        RECT 137.670 111.190 137.930 112.840 ;
        RECT 154.660 112.150 155.540 112.320 ;
        RECT 154.240 111.930 154.410 112.100 ;
        RECT 155.790 111.930 155.960 112.100 ;
        RECT 154.660 111.710 155.540 111.880 ;
        RECT 158.005 112.160 158.885 112.330 ;
        RECT 157.540 111.940 157.710 112.110 ;
        RECT 159.180 111.940 159.350 112.110 ;
        RECT 158.005 111.720 158.885 111.890 ;
        RECT 159.720 111.200 159.980 112.850 ;
        RECT 132.610 110.040 133.490 110.210 ;
        RECT 132.190 109.820 132.360 109.990 ;
        RECT 133.740 109.820 133.910 109.990 ;
        RECT 132.610 109.600 133.490 109.770 ;
        RECT 135.955 110.050 136.835 110.220 ;
        RECT 135.490 109.830 135.660 110.000 ;
        RECT 137.130 109.830 137.300 110.000 ;
        RECT 135.955 109.610 136.835 109.780 ;
        RECT 137.670 109.090 137.930 110.740 ;
        RECT 154.660 110.050 155.540 110.220 ;
        RECT 154.240 109.830 154.410 110.000 ;
        RECT 155.790 109.830 155.960 110.000 ;
        RECT 154.660 109.610 155.540 109.780 ;
        RECT 158.005 110.060 158.885 110.230 ;
        RECT 157.540 109.840 157.710 110.010 ;
        RECT 159.180 109.840 159.350 110.010 ;
        RECT 158.005 109.620 158.885 109.790 ;
        RECT 159.720 109.100 159.980 110.750 ;
        RECT 132.610 107.940 133.490 108.110 ;
        RECT 132.190 107.720 132.360 107.890 ;
        RECT 133.740 107.720 133.910 107.890 ;
        RECT 132.610 107.500 133.490 107.670 ;
        RECT 135.955 107.950 136.835 108.120 ;
        RECT 135.490 107.730 135.660 107.900 ;
        RECT 137.130 107.730 137.300 107.900 ;
        RECT 135.955 107.510 136.835 107.680 ;
        RECT 137.670 106.990 137.930 108.640 ;
        RECT 154.660 107.950 155.540 108.120 ;
        RECT 154.240 107.730 154.410 107.900 ;
        RECT 155.790 107.730 155.960 107.900 ;
        RECT 154.660 107.510 155.540 107.680 ;
        RECT 158.005 107.960 158.885 108.130 ;
        RECT 157.540 107.740 157.710 107.910 ;
        RECT 159.180 107.740 159.350 107.910 ;
        RECT 158.005 107.520 158.885 107.690 ;
        RECT 159.720 107.000 159.980 108.650 ;
        RECT 132.610 105.840 133.490 106.010 ;
        RECT 132.190 105.620 132.360 105.790 ;
        RECT 133.740 105.620 133.910 105.790 ;
        RECT 132.610 105.400 133.490 105.570 ;
        RECT 135.955 105.850 136.835 106.020 ;
        RECT 135.490 105.630 135.660 105.800 ;
        RECT 137.130 105.630 137.300 105.800 ;
        RECT 135.955 105.410 136.835 105.580 ;
        RECT 137.670 104.890 137.930 106.540 ;
        RECT 154.660 105.850 155.540 106.020 ;
        RECT 154.240 105.630 154.410 105.800 ;
        RECT 155.790 105.630 155.960 105.800 ;
        RECT 154.660 105.410 155.540 105.580 ;
        RECT 158.005 105.860 158.885 106.030 ;
        RECT 157.540 105.640 157.710 105.810 ;
        RECT 159.180 105.640 159.350 105.810 ;
        RECT 158.005 105.420 158.885 105.590 ;
        RECT 159.720 104.900 159.980 106.550 ;
        RECT 132.610 103.740 133.490 103.910 ;
        RECT 132.190 103.520 132.360 103.690 ;
        RECT 133.740 103.520 133.910 103.690 ;
        RECT 132.610 103.300 133.490 103.470 ;
        RECT 135.955 103.750 136.835 103.920 ;
        RECT 135.490 103.530 135.660 103.700 ;
        RECT 137.130 103.530 137.300 103.700 ;
        RECT 135.955 103.310 136.835 103.480 ;
        RECT 137.670 102.790 137.930 104.440 ;
        RECT 154.660 103.750 155.540 103.920 ;
        RECT 154.240 103.530 154.410 103.700 ;
        RECT 155.790 103.530 155.960 103.700 ;
        RECT 154.660 103.310 155.540 103.480 ;
        RECT 158.005 103.760 158.885 103.930 ;
        RECT 157.540 103.540 157.710 103.710 ;
        RECT 159.180 103.540 159.350 103.710 ;
        RECT 158.005 103.320 158.885 103.490 ;
        RECT 159.720 102.800 159.980 104.450 ;
        RECT 132.610 101.640 133.490 101.810 ;
        RECT 132.190 101.420 132.360 101.590 ;
        RECT 133.740 101.420 133.910 101.590 ;
        RECT 132.610 101.200 133.490 101.370 ;
        RECT 135.955 101.650 136.835 101.820 ;
        RECT 135.490 101.430 135.660 101.600 ;
        RECT 137.130 101.430 137.300 101.600 ;
        RECT 135.955 101.210 136.835 101.380 ;
        RECT 137.670 100.690 137.930 102.340 ;
        RECT 154.660 101.650 155.540 101.820 ;
        RECT 154.240 101.430 154.410 101.600 ;
        RECT 155.790 101.430 155.960 101.600 ;
        RECT 154.660 101.210 155.540 101.380 ;
        RECT 158.005 101.660 158.885 101.830 ;
        RECT 157.540 101.440 157.710 101.610 ;
        RECT 159.180 101.440 159.350 101.610 ;
        RECT 158.005 101.220 158.885 101.390 ;
        RECT 159.720 100.700 159.980 102.350 ;
        RECT 132.610 99.540 133.490 99.710 ;
        RECT 132.190 99.320 132.360 99.490 ;
        RECT 133.740 99.320 133.910 99.490 ;
        RECT 132.610 99.100 133.490 99.270 ;
        RECT 135.955 99.550 136.835 99.720 ;
        RECT 135.490 99.330 135.660 99.500 ;
        RECT 137.130 99.330 137.300 99.500 ;
        RECT 135.955 99.110 136.835 99.280 ;
        RECT 137.670 98.590 137.930 100.240 ;
        RECT 154.660 99.550 155.540 99.720 ;
        RECT 154.240 99.330 154.410 99.500 ;
        RECT 155.790 99.330 155.960 99.500 ;
        RECT 154.660 99.110 155.540 99.280 ;
        RECT 158.005 99.560 158.885 99.730 ;
        RECT 157.540 99.340 157.710 99.510 ;
        RECT 159.180 99.340 159.350 99.510 ;
        RECT 158.005 99.120 158.885 99.290 ;
        RECT 159.720 98.600 159.980 100.250 ;
        RECT 132.610 97.440 133.490 97.610 ;
        RECT 132.190 97.220 132.360 97.390 ;
        RECT 133.740 97.220 133.910 97.390 ;
        RECT 132.610 97.000 133.490 97.170 ;
        RECT 135.955 97.450 136.835 97.620 ;
        RECT 135.490 97.230 135.660 97.400 ;
        RECT 137.130 97.230 137.300 97.400 ;
        RECT 135.955 97.010 136.835 97.180 ;
        RECT 137.670 96.490 137.930 98.140 ;
        RECT 154.660 97.450 155.540 97.620 ;
        RECT 154.240 97.230 154.410 97.400 ;
        RECT 155.790 97.230 155.960 97.400 ;
        RECT 154.660 97.010 155.540 97.180 ;
        RECT 158.005 97.460 158.885 97.630 ;
        RECT 157.540 97.240 157.710 97.410 ;
        RECT 159.180 97.240 159.350 97.410 ;
        RECT 158.005 97.020 158.885 97.190 ;
        RECT 159.720 96.500 159.980 98.150 ;
        RECT 132.610 95.340 133.490 95.510 ;
        RECT 132.190 95.120 132.360 95.290 ;
        RECT 133.740 95.120 133.910 95.290 ;
        RECT 132.610 94.900 133.490 95.070 ;
        RECT 135.955 95.350 136.835 95.520 ;
        RECT 135.490 95.130 135.660 95.300 ;
        RECT 137.130 95.130 137.300 95.300 ;
        RECT 135.955 94.910 136.835 95.080 ;
        RECT 137.670 94.390 137.930 96.040 ;
        RECT 154.660 95.350 155.540 95.520 ;
        RECT 154.240 95.130 154.410 95.300 ;
        RECT 155.790 95.130 155.960 95.300 ;
        RECT 154.660 94.910 155.540 95.080 ;
        RECT 158.005 95.360 158.885 95.530 ;
        RECT 157.540 95.140 157.710 95.310 ;
        RECT 159.180 95.140 159.350 95.310 ;
        RECT 158.005 94.920 158.885 95.090 ;
        RECT 159.720 94.400 159.980 96.050 ;
        RECT 132.610 93.240 133.490 93.410 ;
        RECT 132.190 93.020 132.360 93.190 ;
        RECT 133.740 93.020 133.910 93.190 ;
        RECT 132.610 92.800 133.490 92.970 ;
        RECT 135.955 93.250 136.835 93.420 ;
        RECT 135.490 93.030 135.660 93.200 ;
        RECT 137.130 93.030 137.300 93.200 ;
        RECT 135.955 92.810 136.835 92.980 ;
        RECT 137.670 92.290 137.930 93.940 ;
        RECT 154.660 93.250 155.540 93.420 ;
        RECT 154.240 93.030 154.410 93.200 ;
        RECT 155.790 93.030 155.960 93.200 ;
        RECT 154.660 92.810 155.540 92.980 ;
        RECT 158.005 93.260 158.885 93.430 ;
        RECT 157.540 93.040 157.710 93.210 ;
        RECT 159.180 93.040 159.350 93.210 ;
        RECT 158.005 92.820 158.885 92.990 ;
        RECT 159.720 92.300 159.980 93.950 ;
        RECT 132.610 91.140 133.490 91.310 ;
        RECT 132.190 90.920 132.360 91.090 ;
        RECT 133.740 90.920 133.910 91.090 ;
        RECT 132.610 90.700 133.490 90.870 ;
        RECT 135.955 91.150 136.835 91.320 ;
        RECT 135.490 90.930 135.660 91.100 ;
        RECT 137.130 90.930 137.300 91.100 ;
        RECT 135.955 90.710 136.835 90.880 ;
        RECT 137.670 90.190 137.930 91.840 ;
        RECT 154.660 91.150 155.540 91.320 ;
        RECT 154.240 90.930 154.410 91.100 ;
        RECT 155.790 90.930 155.960 91.100 ;
        RECT 154.660 90.710 155.540 90.880 ;
        RECT 158.005 91.160 158.885 91.330 ;
        RECT 157.540 90.940 157.710 91.110 ;
        RECT 159.180 90.940 159.350 91.110 ;
        RECT 158.005 90.720 158.885 90.890 ;
        RECT 159.720 90.200 159.980 91.850 ;
        RECT 132.610 89.040 133.490 89.210 ;
        RECT 132.190 88.820 132.360 88.990 ;
        RECT 133.740 88.820 133.910 88.990 ;
        RECT 132.610 88.600 133.490 88.770 ;
        RECT 135.955 89.050 136.835 89.220 ;
        RECT 135.490 88.830 135.660 89.000 ;
        RECT 137.130 88.830 137.300 89.000 ;
        RECT 135.955 88.610 136.835 88.780 ;
        RECT 137.670 88.090 137.930 89.740 ;
        RECT 154.660 89.050 155.540 89.220 ;
        RECT 154.240 88.830 154.410 89.000 ;
        RECT 155.790 88.830 155.960 89.000 ;
        RECT 154.660 88.610 155.540 88.780 ;
        RECT 158.005 89.060 158.885 89.230 ;
        RECT 157.540 88.840 157.710 89.010 ;
        RECT 159.180 88.840 159.350 89.010 ;
        RECT 158.005 88.620 158.885 88.790 ;
        RECT 159.720 88.100 159.980 89.750 ;
        RECT 132.610 86.940 133.490 87.110 ;
        RECT 132.190 86.720 132.360 86.890 ;
        RECT 133.740 86.720 133.910 86.890 ;
        RECT 132.610 86.500 133.490 86.670 ;
        RECT 135.955 86.950 136.835 87.120 ;
        RECT 135.490 86.730 135.660 86.900 ;
        RECT 137.130 86.730 137.300 86.900 ;
        RECT 135.955 86.510 136.835 86.680 ;
        RECT 137.670 85.990 137.930 87.640 ;
        RECT 154.660 86.950 155.540 87.120 ;
        RECT 154.240 86.730 154.410 86.900 ;
        RECT 155.790 86.730 155.960 86.900 ;
        RECT 154.660 86.510 155.540 86.680 ;
        RECT 158.005 86.960 158.885 87.130 ;
        RECT 157.540 86.740 157.710 86.910 ;
        RECT 159.180 86.740 159.350 86.910 ;
        RECT 158.005 86.520 158.885 86.690 ;
        RECT 159.720 86.000 159.980 87.650 ;
        RECT 132.610 84.840 133.490 85.010 ;
        RECT 132.190 84.620 132.360 84.790 ;
        RECT 133.740 84.620 133.910 84.790 ;
        RECT 132.610 84.400 133.490 84.570 ;
        RECT 135.955 84.850 136.835 85.020 ;
        RECT 135.490 84.630 135.660 84.800 ;
        RECT 137.130 84.630 137.300 84.800 ;
        RECT 135.955 84.410 136.835 84.580 ;
        RECT 137.670 83.890 137.930 85.540 ;
        RECT 154.660 84.850 155.540 85.020 ;
        RECT 154.240 84.630 154.410 84.800 ;
        RECT 155.790 84.630 155.960 84.800 ;
        RECT 154.660 84.410 155.540 84.580 ;
        RECT 158.005 84.860 158.885 85.030 ;
        RECT 157.540 84.640 157.710 84.810 ;
        RECT 159.180 84.640 159.350 84.810 ;
        RECT 158.005 84.420 158.885 84.590 ;
        RECT 159.720 83.900 159.980 85.550 ;
        RECT 132.610 82.740 133.490 82.910 ;
        RECT 132.190 82.520 132.360 82.690 ;
        RECT 133.740 82.520 133.910 82.690 ;
        RECT 132.610 82.300 133.490 82.470 ;
        RECT 135.955 82.750 136.835 82.920 ;
        RECT 135.490 82.530 135.660 82.700 ;
        RECT 137.130 82.530 137.300 82.700 ;
        RECT 135.955 82.310 136.835 82.480 ;
        RECT 137.670 81.790 137.930 83.440 ;
        RECT 154.660 82.750 155.540 82.920 ;
        RECT 154.240 82.530 154.410 82.700 ;
        RECT 155.790 82.530 155.960 82.700 ;
        RECT 154.660 82.310 155.540 82.480 ;
        RECT 158.005 82.760 158.885 82.930 ;
        RECT 157.540 82.540 157.710 82.710 ;
        RECT 159.180 82.540 159.350 82.710 ;
        RECT 158.005 82.320 158.885 82.490 ;
        RECT 159.720 81.800 159.980 83.450 ;
        RECT 132.610 80.640 133.490 80.810 ;
        RECT 132.190 80.420 132.360 80.590 ;
        RECT 133.740 80.420 133.910 80.590 ;
        RECT 132.610 80.200 133.490 80.370 ;
        RECT 135.955 80.650 136.835 80.820 ;
        RECT 135.490 80.430 135.660 80.600 ;
        RECT 137.130 80.430 137.300 80.600 ;
        RECT 135.955 80.210 136.835 80.380 ;
        RECT 137.670 79.690 137.930 81.340 ;
        RECT 154.660 80.650 155.540 80.820 ;
        RECT 154.240 80.430 154.410 80.600 ;
        RECT 155.790 80.430 155.960 80.600 ;
        RECT 154.660 80.210 155.540 80.380 ;
        RECT 158.005 80.660 158.885 80.830 ;
        RECT 157.540 80.440 157.710 80.610 ;
        RECT 159.180 80.440 159.350 80.610 ;
        RECT 158.005 80.220 158.885 80.390 ;
        RECT 159.720 79.700 159.980 81.350 ;
        RECT 132.610 78.540 133.490 78.710 ;
        RECT 132.190 78.320 132.360 78.490 ;
        RECT 133.740 78.320 133.910 78.490 ;
        RECT 132.610 78.100 133.490 78.270 ;
        RECT 135.955 78.550 136.835 78.720 ;
        RECT 135.490 78.330 135.660 78.500 ;
        RECT 137.130 78.330 137.300 78.500 ;
        RECT 135.955 78.110 136.835 78.280 ;
        RECT 137.670 77.590 137.930 79.240 ;
        RECT 154.660 78.550 155.540 78.720 ;
        RECT 154.240 78.330 154.410 78.500 ;
        RECT 155.790 78.330 155.960 78.500 ;
        RECT 154.660 78.110 155.540 78.280 ;
        RECT 158.005 78.560 158.885 78.730 ;
        RECT 157.540 78.340 157.710 78.510 ;
        RECT 159.180 78.340 159.350 78.510 ;
        RECT 158.005 78.120 158.885 78.290 ;
        RECT 159.720 77.600 159.980 79.250 ;
        RECT 132.610 76.440 133.490 76.610 ;
        RECT 132.190 76.220 132.360 76.390 ;
        RECT 133.740 76.220 133.910 76.390 ;
        RECT 132.610 76.000 133.490 76.170 ;
        RECT 135.955 76.450 136.835 76.620 ;
        RECT 135.490 76.230 135.660 76.400 ;
        RECT 137.130 76.230 137.300 76.400 ;
        RECT 135.955 76.010 136.835 76.180 ;
        RECT 137.670 75.490 137.930 77.140 ;
        RECT 154.660 76.450 155.540 76.620 ;
        RECT 154.240 76.230 154.410 76.400 ;
        RECT 155.790 76.230 155.960 76.400 ;
        RECT 154.660 76.010 155.540 76.180 ;
        RECT 158.005 76.460 158.885 76.630 ;
        RECT 157.540 76.240 157.710 76.410 ;
        RECT 159.180 76.240 159.350 76.410 ;
        RECT 158.005 76.020 158.885 76.190 ;
        RECT 159.720 75.500 159.980 77.150 ;
        RECT 132.610 74.340 133.490 74.510 ;
        RECT 132.190 74.120 132.360 74.290 ;
        RECT 133.740 74.120 133.910 74.290 ;
        RECT 132.610 73.900 133.490 74.070 ;
        RECT 135.955 74.350 136.835 74.520 ;
        RECT 135.490 74.130 135.660 74.300 ;
        RECT 137.130 74.130 137.300 74.300 ;
        RECT 135.955 73.910 136.835 74.080 ;
        RECT 137.670 73.390 137.930 75.040 ;
        RECT 154.660 74.350 155.540 74.520 ;
        RECT 154.240 74.130 154.410 74.300 ;
        RECT 155.790 74.130 155.960 74.300 ;
        RECT 154.660 73.910 155.540 74.080 ;
        RECT 158.005 74.360 158.885 74.530 ;
        RECT 157.540 74.140 157.710 74.310 ;
        RECT 159.180 74.140 159.350 74.310 ;
        RECT 158.005 73.920 158.885 74.090 ;
        RECT 159.720 73.400 159.980 75.050 ;
        RECT 132.610 72.240 133.490 72.410 ;
        RECT 132.190 72.020 132.360 72.190 ;
        RECT 133.740 72.020 133.910 72.190 ;
        RECT 132.610 71.800 133.490 71.970 ;
        RECT 135.955 72.250 136.835 72.420 ;
        RECT 135.490 72.030 135.660 72.200 ;
        RECT 137.130 72.030 137.300 72.200 ;
        RECT 135.955 71.810 136.835 71.980 ;
        RECT 137.670 71.290 137.930 72.940 ;
        RECT 154.660 72.250 155.540 72.420 ;
        RECT 154.240 72.030 154.410 72.200 ;
        RECT 155.790 72.030 155.960 72.200 ;
        RECT 154.660 71.810 155.540 71.980 ;
        RECT 158.005 72.260 158.885 72.430 ;
        RECT 157.540 72.040 157.710 72.210 ;
        RECT 159.180 72.040 159.350 72.210 ;
        RECT 158.005 71.820 158.885 71.990 ;
        RECT 159.720 71.300 159.980 72.950 ;
        RECT 132.610 70.140 133.490 70.310 ;
        RECT 132.190 69.920 132.360 70.090 ;
        RECT 133.740 69.920 133.910 70.090 ;
        RECT 132.610 69.700 133.490 69.870 ;
        RECT 135.955 70.150 136.835 70.320 ;
        RECT 135.490 69.930 135.660 70.100 ;
        RECT 137.130 69.930 137.300 70.100 ;
        RECT 135.955 69.710 136.835 69.880 ;
        RECT 137.670 69.190 137.930 70.840 ;
        RECT 154.660 70.150 155.540 70.320 ;
        RECT 154.240 69.930 154.410 70.100 ;
        RECT 155.790 69.930 155.960 70.100 ;
        RECT 154.660 69.710 155.540 69.880 ;
        RECT 158.005 70.160 158.885 70.330 ;
        RECT 157.540 69.940 157.710 70.110 ;
        RECT 159.180 69.940 159.350 70.110 ;
        RECT 158.005 69.720 158.885 69.890 ;
        RECT 159.720 69.200 159.980 70.850 ;
        RECT 132.610 68.040 133.490 68.210 ;
        RECT 132.190 67.820 132.360 67.990 ;
        RECT 133.740 67.820 133.910 67.990 ;
        RECT 132.610 67.600 133.490 67.770 ;
        RECT 135.955 68.050 136.835 68.220 ;
        RECT 135.490 67.830 135.660 68.000 ;
        RECT 137.130 67.830 137.300 68.000 ;
        RECT 135.955 67.610 136.835 67.780 ;
        RECT 137.670 67.090 137.930 68.740 ;
        RECT 154.660 68.050 155.540 68.220 ;
        RECT 154.240 67.830 154.410 68.000 ;
        RECT 155.790 67.830 155.960 68.000 ;
        RECT 154.660 67.610 155.540 67.780 ;
        RECT 158.005 68.060 158.885 68.230 ;
        RECT 157.540 67.840 157.710 68.010 ;
        RECT 159.180 67.840 159.350 68.010 ;
        RECT 158.005 67.620 158.885 67.790 ;
        RECT 159.720 67.100 159.980 68.750 ;
        RECT 132.610 65.940 133.490 66.110 ;
        RECT 132.190 65.720 132.360 65.890 ;
        RECT 133.740 65.720 133.910 65.890 ;
        RECT 132.610 65.500 133.490 65.670 ;
        RECT 135.955 65.950 136.835 66.120 ;
        RECT 135.490 65.730 135.660 65.900 ;
        RECT 137.130 65.730 137.300 65.900 ;
        RECT 135.955 65.510 136.835 65.680 ;
        RECT 137.670 64.990 137.930 66.640 ;
        RECT 154.660 65.950 155.540 66.120 ;
        RECT 154.240 65.730 154.410 65.900 ;
        RECT 155.790 65.730 155.960 65.900 ;
        RECT 154.660 65.510 155.540 65.680 ;
        RECT 158.005 65.960 158.885 66.130 ;
        RECT 157.540 65.740 157.710 65.910 ;
        RECT 159.180 65.740 159.350 65.910 ;
        RECT 158.005 65.520 158.885 65.690 ;
        RECT 159.720 65.000 159.980 66.650 ;
        RECT 132.610 63.840 133.490 64.010 ;
        RECT 132.190 63.620 132.360 63.790 ;
        RECT 133.740 63.620 133.910 63.790 ;
        RECT 132.610 63.400 133.490 63.570 ;
        RECT 135.955 63.850 136.835 64.020 ;
        RECT 135.490 63.630 135.660 63.800 ;
        RECT 137.130 63.630 137.300 63.800 ;
        RECT 135.955 63.410 136.835 63.580 ;
        RECT 137.670 62.890 137.930 64.540 ;
        RECT 154.660 63.850 155.540 64.020 ;
        RECT 154.240 63.630 154.410 63.800 ;
        RECT 155.790 63.630 155.960 63.800 ;
        RECT 154.660 63.410 155.540 63.580 ;
        RECT 158.005 63.860 158.885 64.030 ;
        RECT 157.540 63.640 157.710 63.810 ;
        RECT 159.180 63.640 159.350 63.810 ;
        RECT 158.005 63.420 158.885 63.590 ;
        RECT 159.720 62.900 159.980 64.550 ;
        RECT 132.610 61.740 133.490 61.910 ;
        RECT 132.190 61.520 132.360 61.690 ;
        RECT 133.740 61.520 133.910 61.690 ;
        RECT 132.610 61.300 133.490 61.470 ;
        RECT 135.955 61.750 136.835 61.920 ;
        RECT 135.490 61.530 135.660 61.700 ;
        RECT 137.130 61.530 137.300 61.700 ;
        RECT 135.955 61.310 136.835 61.480 ;
        RECT 137.670 60.790 137.930 62.440 ;
        RECT 154.660 61.750 155.540 61.920 ;
        RECT 154.240 61.530 154.410 61.700 ;
        RECT 155.790 61.530 155.960 61.700 ;
        RECT 154.660 61.310 155.540 61.480 ;
        RECT 158.005 61.760 158.885 61.930 ;
        RECT 157.540 61.540 157.710 61.710 ;
        RECT 159.180 61.540 159.350 61.710 ;
        RECT 158.005 61.320 158.885 61.490 ;
        RECT 159.720 60.800 159.980 62.450 ;
        RECT 132.610 59.640 133.490 59.810 ;
        RECT 132.190 59.420 132.360 59.590 ;
        RECT 133.740 59.420 133.910 59.590 ;
        RECT 132.610 59.200 133.490 59.370 ;
        RECT 135.955 59.650 136.835 59.820 ;
        RECT 135.490 59.430 135.660 59.600 ;
        RECT 137.130 59.430 137.300 59.600 ;
        RECT 135.955 59.210 136.835 59.380 ;
        RECT 137.670 58.690 137.930 60.340 ;
        RECT 154.660 59.650 155.540 59.820 ;
        RECT 154.240 59.430 154.410 59.600 ;
        RECT 155.790 59.430 155.960 59.600 ;
        RECT 154.660 59.210 155.540 59.380 ;
        RECT 158.005 59.660 158.885 59.830 ;
        RECT 157.540 59.440 157.710 59.610 ;
        RECT 159.180 59.440 159.350 59.610 ;
        RECT 158.005 59.220 158.885 59.390 ;
        RECT 159.720 58.700 159.980 60.350 ;
        RECT 132.610 57.540 133.490 57.710 ;
        RECT 132.190 57.320 132.360 57.490 ;
        RECT 133.740 57.320 133.910 57.490 ;
        RECT 132.610 57.100 133.490 57.270 ;
        RECT 135.955 57.550 136.835 57.720 ;
        RECT 135.490 57.330 135.660 57.500 ;
        RECT 137.130 57.330 137.300 57.500 ;
        RECT 135.955 57.110 136.835 57.280 ;
        RECT 137.670 56.590 137.930 58.240 ;
        RECT 154.660 57.550 155.540 57.720 ;
        RECT 154.240 57.330 154.410 57.500 ;
        RECT 155.790 57.330 155.960 57.500 ;
        RECT 154.660 57.110 155.540 57.280 ;
        RECT 158.005 57.560 158.885 57.730 ;
        RECT 157.540 57.340 157.710 57.510 ;
        RECT 159.180 57.340 159.350 57.510 ;
        RECT 158.005 57.120 158.885 57.290 ;
        RECT 159.720 56.600 159.980 58.250 ;
        RECT 132.610 55.440 133.490 55.610 ;
        RECT 132.190 55.220 132.360 55.390 ;
        RECT 133.740 55.220 133.910 55.390 ;
        RECT 132.610 55.000 133.490 55.170 ;
        RECT 135.955 55.450 136.835 55.620 ;
        RECT 135.490 55.230 135.660 55.400 ;
        RECT 137.130 55.230 137.300 55.400 ;
        RECT 135.955 55.010 136.835 55.180 ;
        RECT 137.670 54.490 137.930 56.140 ;
        RECT 154.660 55.450 155.540 55.620 ;
        RECT 154.240 55.230 154.410 55.400 ;
        RECT 155.790 55.230 155.960 55.400 ;
        RECT 154.660 55.010 155.540 55.180 ;
        RECT 158.005 55.460 158.885 55.630 ;
        RECT 157.540 55.240 157.710 55.410 ;
        RECT 159.180 55.240 159.350 55.410 ;
        RECT 158.005 55.020 158.885 55.190 ;
        RECT 159.720 54.500 159.980 56.150 ;
        RECT 132.610 53.340 133.490 53.510 ;
        RECT 132.190 53.120 132.360 53.290 ;
        RECT 133.740 53.120 133.910 53.290 ;
        RECT 132.610 52.900 133.490 53.070 ;
        RECT 135.955 53.350 136.835 53.520 ;
        RECT 135.490 53.130 135.660 53.300 ;
        RECT 137.130 53.130 137.300 53.300 ;
        RECT 135.955 52.910 136.835 53.080 ;
        RECT 137.670 52.390 137.930 54.040 ;
        RECT 154.660 53.350 155.540 53.520 ;
        RECT 154.240 53.130 154.410 53.300 ;
        RECT 155.790 53.130 155.960 53.300 ;
        RECT 154.660 52.910 155.540 53.080 ;
        RECT 158.005 53.360 158.885 53.530 ;
        RECT 157.540 53.140 157.710 53.310 ;
        RECT 159.180 53.140 159.350 53.310 ;
        RECT 158.005 52.920 158.885 53.090 ;
        RECT 159.720 52.400 159.980 54.050 ;
        RECT 132.610 51.240 133.490 51.410 ;
        RECT 132.190 51.020 132.360 51.190 ;
        RECT 133.740 51.020 133.910 51.190 ;
        RECT 132.610 50.800 133.490 50.970 ;
        RECT 135.955 51.250 136.835 51.420 ;
        RECT 135.490 51.030 135.660 51.200 ;
        RECT 137.130 51.030 137.300 51.200 ;
        RECT 135.955 50.810 136.835 50.980 ;
        RECT 137.670 50.290 137.930 51.940 ;
        RECT 154.660 51.250 155.540 51.420 ;
        RECT 154.240 51.030 154.410 51.200 ;
        RECT 155.790 51.030 155.960 51.200 ;
        RECT 154.660 50.810 155.540 50.980 ;
        RECT 158.005 51.260 158.885 51.430 ;
        RECT 157.540 51.040 157.710 51.210 ;
        RECT 159.180 51.040 159.350 51.210 ;
        RECT 158.005 50.820 158.885 50.990 ;
        RECT 159.720 50.300 159.980 51.950 ;
        RECT 132.610 49.140 133.490 49.310 ;
        RECT 132.190 48.920 132.360 49.090 ;
        RECT 133.740 48.920 133.910 49.090 ;
        RECT 132.610 48.700 133.490 48.870 ;
        RECT 135.955 49.150 136.835 49.320 ;
        RECT 135.490 48.930 135.660 49.100 ;
        RECT 137.130 48.930 137.300 49.100 ;
        RECT 135.955 48.710 136.835 48.880 ;
        RECT 137.670 48.190 137.930 49.840 ;
        RECT 154.660 49.150 155.540 49.320 ;
        RECT 154.240 48.930 154.410 49.100 ;
        RECT 155.790 48.930 155.960 49.100 ;
        RECT 154.660 48.710 155.540 48.880 ;
        RECT 158.005 49.160 158.885 49.330 ;
        RECT 157.540 48.940 157.710 49.110 ;
        RECT 159.180 48.940 159.350 49.110 ;
        RECT 158.005 48.720 158.885 48.890 ;
        RECT 159.720 48.200 159.980 49.850 ;
        RECT 132.610 47.040 133.490 47.210 ;
        RECT 132.190 46.820 132.360 46.990 ;
        RECT 133.740 46.820 133.910 46.990 ;
        RECT 132.610 46.600 133.490 46.770 ;
        RECT 135.955 47.050 136.835 47.220 ;
        RECT 135.490 46.830 135.660 47.000 ;
        RECT 137.130 46.830 137.300 47.000 ;
        RECT 135.955 46.610 136.835 46.780 ;
        RECT 137.670 46.090 137.930 47.740 ;
        RECT 154.660 47.050 155.540 47.220 ;
        RECT 154.240 46.830 154.410 47.000 ;
        RECT 155.790 46.830 155.960 47.000 ;
        RECT 154.660 46.610 155.540 46.780 ;
        RECT 158.005 47.060 158.885 47.230 ;
        RECT 157.540 46.840 157.710 47.010 ;
        RECT 159.180 46.840 159.350 47.010 ;
        RECT 158.005 46.620 158.885 46.790 ;
        RECT 159.720 46.100 159.980 47.750 ;
        RECT 132.610 44.940 133.490 45.110 ;
        RECT 132.190 44.720 132.360 44.890 ;
        RECT 133.740 44.720 133.910 44.890 ;
        RECT 132.610 44.500 133.490 44.670 ;
        RECT 135.955 44.950 136.835 45.120 ;
        RECT 135.490 44.730 135.660 44.900 ;
        RECT 137.130 44.730 137.300 44.900 ;
        RECT 135.955 44.510 136.835 44.680 ;
        RECT 137.670 43.990 137.930 45.640 ;
        RECT 154.660 44.950 155.540 45.120 ;
        RECT 154.240 44.730 154.410 44.900 ;
        RECT 155.790 44.730 155.960 44.900 ;
        RECT 154.660 44.510 155.540 44.680 ;
        RECT 158.005 44.960 158.885 45.130 ;
        RECT 157.540 44.740 157.710 44.910 ;
        RECT 159.180 44.740 159.350 44.910 ;
        RECT 158.005 44.520 158.885 44.690 ;
        RECT 159.720 44.000 159.980 45.650 ;
        RECT 132.610 42.840 133.490 43.010 ;
        RECT 132.190 42.620 132.360 42.790 ;
        RECT 133.740 42.620 133.910 42.790 ;
        RECT 132.610 42.400 133.490 42.570 ;
        RECT 135.955 42.850 136.835 43.020 ;
        RECT 135.490 42.630 135.660 42.800 ;
        RECT 137.130 42.630 137.300 42.800 ;
        RECT 135.955 42.410 136.835 42.580 ;
        RECT 137.670 41.890 137.930 43.540 ;
        RECT 154.660 42.850 155.540 43.020 ;
        RECT 154.240 42.630 154.410 42.800 ;
        RECT 155.790 42.630 155.960 42.800 ;
        RECT 154.660 42.410 155.540 42.580 ;
        RECT 158.005 42.860 158.885 43.030 ;
        RECT 157.540 42.640 157.710 42.810 ;
        RECT 159.180 42.640 159.350 42.810 ;
        RECT 158.005 42.420 158.885 42.590 ;
        RECT 159.720 41.900 159.980 43.550 ;
        RECT 132.610 40.740 133.490 40.910 ;
        RECT 132.190 40.520 132.360 40.690 ;
        RECT 133.740 40.520 133.910 40.690 ;
        RECT 132.610 40.300 133.490 40.470 ;
        RECT 135.955 40.750 136.835 40.920 ;
        RECT 135.490 40.530 135.660 40.700 ;
        RECT 137.130 40.530 137.300 40.700 ;
        RECT 135.955 40.310 136.835 40.480 ;
        RECT 137.670 39.790 137.930 41.440 ;
        RECT 154.660 40.750 155.540 40.920 ;
        RECT 154.240 40.530 154.410 40.700 ;
        RECT 155.790 40.530 155.960 40.700 ;
        RECT 154.660 40.310 155.540 40.480 ;
        RECT 158.005 40.760 158.885 40.930 ;
        RECT 157.540 40.540 157.710 40.710 ;
        RECT 159.180 40.540 159.350 40.710 ;
        RECT 158.005 40.320 158.885 40.490 ;
        RECT 159.720 39.800 159.980 41.450 ;
        RECT 132.610 38.640 133.490 38.810 ;
        RECT 132.190 38.420 132.360 38.590 ;
        RECT 133.740 38.420 133.910 38.590 ;
        RECT 132.610 38.200 133.490 38.370 ;
        RECT 135.955 38.650 136.835 38.820 ;
        RECT 135.490 38.430 135.660 38.600 ;
        RECT 137.130 38.430 137.300 38.600 ;
        RECT 135.955 38.210 136.835 38.380 ;
        RECT 137.670 37.690 137.930 39.340 ;
        RECT 154.660 38.650 155.540 38.820 ;
        RECT 154.240 38.430 154.410 38.600 ;
        RECT 155.790 38.430 155.960 38.600 ;
        RECT 154.660 38.210 155.540 38.380 ;
        RECT 158.005 38.660 158.885 38.830 ;
        RECT 157.540 38.440 157.710 38.610 ;
        RECT 159.180 38.440 159.350 38.610 ;
        RECT 158.005 38.220 158.885 38.390 ;
        RECT 159.720 37.700 159.980 39.350 ;
        RECT 132.610 36.540 133.490 36.710 ;
        RECT 132.190 36.320 132.360 36.490 ;
        RECT 133.740 36.320 133.910 36.490 ;
        RECT 132.610 36.100 133.490 36.270 ;
        RECT 135.955 36.550 136.835 36.720 ;
        RECT 135.490 36.330 135.660 36.500 ;
        RECT 137.130 36.330 137.300 36.500 ;
        RECT 135.955 36.110 136.835 36.280 ;
        RECT 137.670 35.590 137.930 37.240 ;
        RECT 154.660 36.550 155.540 36.720 ;
        RECT 154.240 36.330 154.410 36.500 ;
        RECT 155.790 36.330 155.960 36.500 ;
        RECT 154.660 36.110 155.540 36.280 ;
        RECT 158.005 36.560 158.885 36.730 ;
        RECT 157.540 36.340 157.710 36.510 ;
        RECT 159.180 36.340 159.350 36.510 ;
        RECT 158.005 36.120 158.885 36.290 ;
        RECT 159.720 35.600 159.980 37.250 ;
        RECT 132.610 34.440 133.490 34.610 ;
        RECT 132.190 34.220 132.360 34.390 ;
        RECT 133.740 34.220 133.910 34.390 ;
        RECT 132.610 34.000 133.490 34.170 ;
        RECT 135.955 34.450 136.835 34.620 ;
        RECT 135.490 34.230 135.660 34.400 ;
        RECT 137.130 34.230 137.300 34.400 ;
        RECT 135.955 34.010 136.835 34.180 ;
        RECT 137.670 33.490 137.930 35.140 ;
        RECT 154.660 34.450 155.540 34.620 ;
        RECT 154.240 34.230 154.410 34.400 ;
        RECT 155.790 34.230 155.960 34.400 ;
        RECT 154.660 34.010 155.540 34.180 ;
        RECT 158.005 34.460 158.885 34.630 ;
        RECT 157.540 34.240 157.710 34.410 ;
        RECT 159.180 34.240 159.350 34.410 ;
        RECT 158.005 34.020 158.885 34.190 ;
        RECT 159.720 33.500 159.980 35.150 ;
        RECT 132.610 32.340 133.490 32.510 ;
        RECT 132.190 32.120 132.360 32.290 ;
        RECT 133.740 32.120 133.910 32.290 ;
        RECT 132.610 31.900 133.490 32.070 ;
        RECT 135.955 32.350 136.835 32.520 ;
        RECT 135.490 32.130 135.660 32.300 ;
        RECT 137.130 32.130 137.300 32.300 ;
        RECT 135.955 31.910 136.835 32.080 ;
        RECT 137.670 31.390 137.930 33.040 ;
        RECT 154.660 32.350 155.540 32.520 ;
        RECT 154.240 32.130 154.410 32.300 ;
        RECT 155.790 32.130 155.960 32.300 ;
        RECT 154.660 31.910 155.540 32.080 ;
        RECT 158.005 32.360 158.885 32.530 ;
        RECT 157.540 32.140 157.710 32.310 ;
        RECT 159.180 32.140 159.350 32.310 ;
        RECT 158.005 31.920 158.885 32.090 ;
        RECT 159.720 31.400 159.980 33.050 ;
        RECT 132.610 30.240 133.490 30.410 ;
        RECT 132.190 30.020 132.360 30.190 ;
        RECT 133.740 30.020 133.910 30.190 ;
        RECT 132.610 29.800 133.490 29.970 ;
        RECT 135.955 30.250 136.835 30.420 ;
        RECT 135.490 30.030 135.660 30.200 ;
        RECT 137.130 30.030 137.300 30.200 ;
        RECT 135.955 29.810 136.835 29.980 ;
        RECT 137.670 29.290 137.930 30.940 ;
        RECT 154.660 30.250 155.540 30.420 ;
        RECT 154.240 30.030 154.410 30.200 ;
        RECT 155.790 30.030 155.960 30.200 ;
        RECT 154.660 29.810 155.540 29.980 ;
        RECT 158.005 30.260 158.885 30.430 ;
        RECT 157.540 30.040 157.710 30.210 ;
        RECT 159.180 30.040 159.350 30.210 ;
        RECT 158.005 29.820 158.885 29.990 ;
        RECT 159.720 29.300 159.980 30.950 ;
        RECT 132.610 28.140 133.490 28.310 ;
        RECT 132.190 27.920 132.360 28.090 ;
        RECT 133.740 27.920 133.910 28.090 ;
        RECT 132.610 27.700 133.490 27.870 ;
        RECT 135.955 28.150 136.835 28.320 ;
        RECT 135.490 27.930 135.660 28.100 ;
        RECT 137.130 27.930 137.300 28.100 ;
        RECT 135.955 27.710 136.835 27.880 ;
        RECT 137.670 27.190 137.930 28.840 ;
        RECT 154.660 28.150 155.540 28.320 ;
        RECT 154.240 27.930 154.410 28.100 ;
        RECT 155.790 27.930 155.960 28.100 ;
        RECT 154.660 27.710 155.540 27.880 ;
        RECT 158.005 28.160 158.885 28.330 ;
        RECT 157.540 27.940 157.710 28.110 ;
        RECT 159.180 27.940 159.350 28.110 ;
        RECT 158.005 27.720 158.885 27.890 ;
        RECT 159.720 27.200 159.980 28.850 ;
        RECT 132.610 26.040 133.490 26.210 ;
        RECT 132.190 25.820 132.360 25.990 ;
        RECT 133.740 25.820 133.910 25.990 ;
        RECT 132.610 25.600 133.490 25.770 ;
        RECT 135.955 26.050 136.835 26.220 ;
        RECT 135.490 25.830 135.660 26.000 ;
        RECT 137.130 25.830 137.300 26.000 ;
        RECT 135.955 25.610 136.835 25.780 ;
        RECT 137.670 25.090 137.930 26.740 ;
        RECT 154.660 26.050 155.540 26.220 ;
        RECT 154.240 25.830 154.410 26.000 ;
        RECT 155.790 25.830 155.960 26.000 ;
        RECT 154.660 25.610 155.540 25.780 ;
        RECT 158.005 26.060 158.885 26.230 ;
        RECT 157.540 25.840 157.710 26.010 ;
        RECT 159.180 25.840 159.350 26.010 ;
        RECT 158.005 25.620 158.885 25.790 ;
        RECT 159.720 25.100 159.980 26.750 ;
        RECT 132.610 23.940 133.490 24.110 ;
        RECT 132.190 23.720 132.360 23.890 ;
        RECT 133.740 23.720 133.910 23.890 ;
        RECT 132.610 23.500 133.490 23.670 ;
        RECT 135.955 23.950 136.835 24.120 ;
        RECT 135.490 23.730 135.660 23.900 ;
        RECT 137.130 23.730 137.300 23.900 ;
        RECT 135.955 23.510 136.835 23.680 ;
        RECT 137.670 22.990 137.930 24.640 ;
        RECT 154.660 23.950 155.540 24.120 ;
        RECT 154.240 23.730 154.410 23.900 ;
        RECT 155.790 23.730 155.960 23.900 ;
        RECT 154.660 23.510 155.540 23.680 ;
        RECT 158.005 23.960 158.885 24.130 ;
        RECT 157.540 23.740 157.710 23.910 ;
        RECT 159.180 23.740 159.350 23.910 ;
        RECT 158.005 23.520 158.885 23.690 ;
        RECT 159.720 23.000 159.980 24.650 ;
        RECT 132.610 21.840 133.490 22.010 ;
        RECT 132.190 21.620 132.360 21.790 ;
        RECT 133.740 21.620 133.910 21.790 ;
        RECT 132.610 21.400 133.490 21.570 ;
        RECT 135.955 21.850 136.835 22.020 ;
        RECT 135.490 21.630 135.660 21.800 ;
        RECT 137.130 21.630 137.300 21.800 ;
        RECT 135.955 21.410 136.835 21.580 ;
        RECT 137.670 20.890 137.930 22.540 ;
        RECT 154.660 21.850 155.540 22.020 ;
        RECT 154.240 21.630 154.410 21.800 ;
        RECT 155.790 21.630 155.960 21.800 ;
        RECT 154.660 21.410 155.540 21.580 ;
        RECT 158.005 21.860 158.885 22.030 ;
        RECT 157.540 21.640 157.710 21.810 ;
        RECT 159.180 21.640 159.350 21.810 ;
        RECT 158.005 21.420 158.885 21.590 ;
        RECT 159.720 20.900 159.980 22.550 ;
        RECT 132.610 19.740 133.490 19.910 ;
        RECT 132.190 19.520 132.360 19.690 ;
        RECT 133.740 19.520 133.910 19.690 ;
        RECT 132.610 19.300 133.490 19.470 ;
        RECT 135.955 19.750 136.835 19.920 ;
        RECT 135.490 19.530 135.660 19.700 ;
        RECT 137.130 19.530 137.300 19.700 ;
        RECT 135.955 19.310 136.835 19.480 ;
        RECT 137.670 18.790 137.930 20.440 ;
        RECT 154.660 19.750 155.540 19.920 ;
        RECT 154.240 19.530 154.410 19.700 ;
        RECT 155.790 19.530 155.960 19.700 ;
        RECT 154.660 19.310 155.540 19.480 ;
        RECT 158.005 19.760 158.885 19.930 ;
        RECT 157.540 19.540 157.710 19.710 ;
        RECT 159.180 19.540 159.350 19.710 ;
        RECT 158.005 19.320 158.885 19.490 ;
        RECT 159.720 18.800 159.980 20.450 ;
        RECT 132.610 17.640 133.490 17.810 ;
        RECT 132.190 17.420 132.360 17.590 ;
        RECT 133.740 17.420 133.910 17.590 ;
        RECT 132.610 17.200 133.490 17.370 ;
        RECT 135.955 17.650 136.835 17.820 ;
        RECT 135.490 17.430 135.660 17.600 ;
        RECT 137.130 17.430 137.300 17.600 ;
        RECT 135.955 17.210 136.835 17.380 ;
        RECT 137.670 16.690 137.930 18.340 ;
        RECT 154.660 17.650 155.540 17.820 ;
        RECT 154.240 17.430 154.410 17.600 ;
        RECT 155.790 17.430 155.960 17.600 ;
        RECT 154.660 17.210 155.540 17.380 ;
        RECT 158.005 17.660 158.885 17.830 ;
        RECT 157.540 17.440 157.710 17.610 ;
        RECT 159.180 17.440 159.350 17.610 ;
        RECT 158.005 17.220 158.885 17.390 ;
        RECT 159.720 16.700 159.980 18.350 ;
        RECT 132.610 15.540 133.490 15.710 ;
        RECT 132.190 15.320 132.360 15.490 ;
        RECT 133.740 15.320 133.910 15.490 ;
        RECT 132.610 15.100 133.490 15.270 ;
        RECT 135.955 15.550 136.835 15.720 ;
        RECT 135.490 15.330 135.660 15.500 ;
        RECT 137.130 15.330 137.300 15.500 ;
        RECT 135.955 15.110 136.835 15.280 ;
        RECT 137.670 14.590 137.930 16.240 ;
        RECT 154.660 15.550 155.540 15.720 ;
        RECT 154.240 15.330 154.410 15.500 ;
        RECT 155.790 15.330 155.960 15.500 ;
        RECT 154.660 15.110 155.540 15.280 ;
        RECT 158.005 15.560 158.885 15.730 ;
        RECT 157.540 15.340 157.710 15.510 ;
        RECT 159.180 15.340 159.350 15.510 ;
        RECT 158.005 15.120 158.885 15.290 ;
        RECT 159.720 14.600 159.980 16.250 ;
        RECT 132.610 13.440 133.490 13.610 ;
        RECT 132.190 13.220 132.360 13.390 ;
        RECT 133.740 13.220 133.910 13.390 ;
        RECT 132.610 13.000 133.490 13.170 ;
        RECT 135.955 13.450 136.835 13.620 ;
        RECT 135.490 13.230 135.660 13.400 ;
        RECT 137.130 13.230 137.300 13.400 ;
        RECT 135.955 13.010 136.835 13.180 ;
        RECT 137.670 12.490 137.930 14.140 ;
        RECT 154.660 13.450 155.540 13.620 ;
        RECT 154.240 13.230 154.410 13.400 ;
        RECT 155.790 13.230 155.960 13.400 ;
        RECT 154.660 13.010 155.540 13.180 ;
        RECT 158.005 13.460 158.885 13.630 ;
        RECT 157.540 13.240 157.710 13.410 ;
        RECT 159.180 13.240 159.350 13.410 ;
        RECT 158.005 13.020 158.885 13.190 ;
        RECT 159.720 12.500 159.980 14.150 ;
        RECT 132.610 11.340 133.490 11.510 ;
        RECT 132.190 11.120 132.360 11.290 ;
        RECT 133.740 11.120 133.910 11.290 ;
        RECT 132.610 10.900 133.490 11.070 ;
        RECT 135.955 11.350 136.835 11.520 ;
        RECT 135.490 11.130 135.660 11.300 ;
        RECT 137.130 11.130 137.300 11.300 ;
        RECT 135.955 10.910 136.835 11.080 ;
        RECT 137.670 10.390 137.930 12.040 ;
        RECT 154.660 11.350 155.540 11.520 ;
        RECT 154.240 11.130 154.410 11.300 ;
        RECT 155.790 11.130 155.960 11.300 ;
        RECT 154.660 10.910 155.540 11.080 ;
        RECT 158.005 11.360 158.885 11.530 ;
        RECT 157.540 11.140 157.710 11.310 ;
        RECT 159.180 11.140 159.350 11.310 ;
        RECT 158.005 10.920 158.885 11.090 ;
        RECT 159.720 10.400 159.980 12.050 ;
        RECT 132.610 9.240 133.490 9.410 ;
        RECT 132.190 9.020 132.360 9.190 ;
        RECT 133.740 9.020 133.910 9.190 ;
        RECT 132.610 8.800 133.490 8.970 ;
        RECT 135.955 9.250 136.835 9.420 ;
        RECT 135.490 9.030 135.660 9.200 ;
        RECT 137.130 9.030 137.300 9.200 ;
        RECT 135.955 8.810 136.835 8.980 ;
        RECT 137.670 8.290 137.930 9.940 ;
        RECT 154.660 9.250 155.540 9.420 ;
        RECT 154.240 9.030 154.410 9.200 ;
        RECT 155.790 9.030 155.960 9.200 ;
        RECT 154.660 8.810 155.540 8.980 ;
        RECT 158.005 9.260 158.885 9.430 ;
        RECT 157.540 9.040 157.710 9.210 ;
        RECT 159.180 9.040 159.350 9.210 ;
        RECT 158.005 8.820 158.885 8.990 ;
        RECT 159.720 8.300 159.980 9.950 ;
        RECT 132.610 7.140 133.490 7.310 ;
        RECT 132.190 6.920 132.360 7.090 ;
        RECT 133.740 6.920 133.910 7.090 ;
        RECT 132.610 6.700 133.490 6.870 ;
        RECT 135.955 7.150 136.835 7.320 ;
        RECT 135.490 6.930 135.660 7.100 ;
        RECT 137.130 6.930 137.300 7.100 ;
        RECT 135.955 6.710 136.835 6.880 ;
        RECT 137.670 6.190 137.930 7.840 ;
        RECT 154.660 7.150 155.540 7.320 ;
        RECT 154.240 6.930 154.410 7.100 ;
        RECT 155.790 6.930 155.960 7.100 ;
        RECT 154.660 6.710 155.540 6.880 ;
        RECT 158.005 7.160 158.885 7.330 ;
        RECT 157.540 6.940 157.710 7.110 ;
        RECT 159.180 6.940 159.350 7.110 ;
        RECT 158.005 6.720 158.885 6.890 ;
        RECT 159.720 6.200 159.980 7.850 ;
        RECT 132.610 5.040 133.490 5.210 ;
        RECT 132.190 4.820 132.360 4.990 ;
        RECT 133.740 4.820 133.910 4.990 ;
        RECT 132.610 4.600 133.490 4.770 ;
        RECT 135.955 5.050 136.835 5.220 ;
        RECT 135.490 4.830 135.660 5.000 ;
        RECT 137.130 4.830 137.300 5.000 ;
        RECT 135.955 4.610 136.835 4.780 ;
        RECT 137.670 4.090 137.930 5.740 ;
        RECT 154.660 5.050 155.540 5.220 ;
        RECT 154.240 4.830 154.410 5.000 ;
        RECT 155.790 4.830 155.960 5.000 ;
        RECT 154.660 4.610 155.540 4.780 ;
        RECT 158.005 5.060 158.885 5.230 ;
        RECT 157.540 4.840 157.710 5.010 ;
        RECT 159.180 4.840 159.350 5.010 ;
        RECT 158.005 4.620 158.885 4.790 ;
        RECT 159.720 4.100 159.980 5.750 ;
        RECT 132.610 2.940 133.490 3.110 ;
        RECT 132.190 2.720 132.360 2.890 ;
        RECT 133.740 2.720 133.910 2.890 ;
        RECT 132.610 2.500 133.490 2.670 ;
        RECT 135.955 2.950 136.835 3.120 ;
        RECT 135.490 2.730 135.660 2.900 ;
        RECT 137.130 2.730 137.300 2.900 ;
        RECT 135.955 2.510 136.835 2.680 ;
        RECT 137.670 1.990 137.930 3.640 ;
        RECT 154.660 2.950 155.540 3.120 ;
        RECT 154.240 2.730 154.410 2.900 ;
        RECT 155.790 2.730 155.960 2.900 ;
        RECT 154.660 2.510 155.540 2.680 ;
        RECT 158.005 2.960 158.885 3.130 ;
        RECT 157.540 2.740 157.710 2.910 ;
        RECT 159.180 2.740 159.350 2.910 ;
        RECT 158.005 2.520 158.885 2.690 ;
        RECT 159.720 2.000 159.980 3.650 ;
      LAYER met1 ;
        RECT 13.740 213.930 19.920 215.050 ;
        RECT 13.740 213.910 114.560 213.930 ;
        RECT 13.740 213.040 160.050 213.910 ;
        RECT 13.740 212.960 114.560 213.040 ;
        RECT 13.740 211.680 19.920 212.960 ;
        RECT 131.250 211.870 131.970 212.720 ;
        RECT 131.490 211.520 131.860 211.870 ;
        RECT 131.490 211.250 133.550 211.520 ;
        RECT 131.490 209.420 131.860 211.250 ;
        RECT 132.110 210.790 132.370 210.820 ;
        RECT 132.110 210.500 132.390 210.790 ;
        RECT 132.550 210.700 133.550 211.250 ;
        RECT 134.420 210.820 135.150 211.690 ;
        RECT 137.640 211.590 137.990 213.040 ;
        RECT 154.050 213.030 154.320 213.040 ;
        RECT 153.170 212.010 154.300 212.650 ;
        RECT 159.700 212.460 160.050 213.040 ;
        RECT 159.690 212.420 160.050 212.460 ;
        RECT 135.870 211.320 137.990 211.590 ;
        RECT 132.550 210.530 133.550 210.540 ;
        RECT 132.110 210.480 132.370 210.500 ;
        RECT 132.540 210.320 133.550 210.530 ;
        RECT 133.690 210.490 135.720 210.820 ;
        RECT 135.880 210.790 136.910 211.320 ;
        RECT 135.895 210.760 136.895 210.790 ;
        RECT 135.895 210.530 136.895 210.550 ;
        RECT 132.540 210.230 133.690 210.320 ;
        RECT 135.870 210.230 136.910 210.530 ;
        RECT 137.070 210.490 137.390 210.820 ;
        RECT 132.540 210.090 136.910 210.230 ;
        RECT 132.540 210.070 135.920 210.090 ;
        RECT 131.490 209.150 133.550 209.420 ;
        RECT 131.490 207.320 131.860 209.150 ;
        RECT 132.110 208.690 132.370 208.720 ;
        RECT 132.110 208.400 132.390 208.690 ;
        RECT 132.550 208.600 133.550 209.150 ;
        RECT 134.420 208.720 135.150 210.070 ;
        RECT 137.640 209.490 137.990 211.320 ;
        RECT 135.870 209.220 137.990 209.490 ;
        RECT 132.550 208.430 133.550 208.440 ;
        RECT 132.110 208.380 132.370 208.400 ;
        RECT 132.540 208.220 133.550 208.430 ;
        RECT 133.690 208.390 135.720 208.720 ;
        RECT 135.880 208.690 136.910 209.220 ;
        RECT 135.895 208.660 136.895 208.690 ;
        RECT 135.895 208.430 136.895 208.450 ;
        RECT 132.540 208.130 133.690 208.220 ;
        RECT 135.870 208.130 136.910 208.430 ;
        RECT 137.070 208.390 137.390 208.720 ;
        RECT 132.540 207.990 136.910 208.130 ;
        RECT 132.540 207.970 135.920 207.990 ;
        RECT 131.490 207.050 133.550 207.320 ;
        RECT 131.490 205.220 131.860 207.050 ;
        RECT 132.110 206.590 132.370 206.620 ;
        RECT 132.110 206.300 132.390 206.590 ;
        RECT 132.550 206.500 133.550 207.050 ;
        RECT 134.420 206.620 135.150 207.970 ;
        RECT 137.640 207.390 137.990 209.220 ;
        RECT 135.870 207.120 137.990 207.390 ;
        RECT 132.550 206.330 133.550 206.340 ;
        RECT 132.110 206.280 132.370 206.300 ;
        RECT 132.540 206.120 133.550 206.330 ;
        RECT 133.690 206.290 135.720 206.620 ;
        RECT 135.880 206.590 136.910 207.120 ;
        RECT 135.895 206.560 136.895 206.590 ;
        RECT 135.895 206.330 136.895 206.350 ;
        RECT 132.540 206.030 133.690 206.120 ;
        RECT 135.870 206.030 136.910 206.330 ;
        RECT 137.070 206.290 137.390 206.620 ;
        RECT 132.540 205.890 136.910 206.030 ;
        RECT 132.540 205.870 135.920 205.890 ;
        RECT 131.490 204.950 133.550 205.220 ;
        RECT 131.490 203.130 131.860 204.950 ;
        RECT 132.110 204.490 132.370 204.520 ;
        RECT 132.110 204.200 132.390 204.490 ;
        RECT 132.550 204.400 133.550 204.950 ;
        RECT 134.420 204.520 135.150 205.870 ;
        RECT 137.640 205.290 137.990 207.120 ;
        RECT 135.870 205.020 137.990 205.290 ;
        RECT 132.550 204.230 133.550 204.240 ;
        RECT 132.110 204.180 132.370 204.200 ;
        RECT 132.540 204.020 133.550 204.230 ;
        RECT 133.690 204.190 135.720 204.520 ;
        RECT 135.880 204.490 136.910 205.020 ;
        RECT 135.895 204.460 136.895 204.490 ;
        RECT 135.895 204.230 136.895 204.250 ;
        RECT 132.540 203.930 133.690 204.020 ;
        RECT 135.870 203.930 136.910 204.230 ;
        RECT 137.070 204.190 137.390 204.520 ;
        RECT 132.540 203.790 136.910 203.930 ;
        RECT 132.540 203.770 135.920 203.790 ;
        RECT 131.490 202.860 133.550 203.130 ;
        RECT 131.490 201.030 131.860 202.860 ;
        RECT 132.110 202.400 132.370 202.430 ;
        RECT 132.110 202.110 132.390 202.400 ;
        RECT 132.550 202.310 133.550 202.860 ;
        RECT 134.420 202.430 135.150 203.770 ;
        RECT 137.640 203.200 137.990 205.020 ;
        RECT 135.870 202.930 137.990 203.200 ;
        RECT 132.550 202.140 133.550 202.150 ;
        RECT 132.110 202.090 132.370 202.110 ;
        RECT 132.540 201.930 133.550 202.140 ;
        RECT 133.690 202.100 135.720 202.430 ;
        RECT 135.880 202.400 136.910 202.930 ;
        RECT 135.895 202.370 136.895 202.400 ;
        RECT 135.895 202.140 136.895 202.160 ;
        RECT 132.540 201.840 133.690 201.930 ;
        RECT 135.870 201.840 136.910 202.140 ;
        RECT 137.070 202.100 137.390 202.430 ;
        RECT 132.540 201.700 136.910 201.840 ;
        RECT 132.540 201.680 135.920 201.700 ;
        RECT 131.490 200.760 133.550 201.030 ;
        RECT 131.490 198.940 131.860 200.760 ;
        RECT 132.110 200.300 132.370 200.330 ;
        RECT 132.110 200.010 132.390 200.300 ;
        RECT 132.550 200.210 133.550 200.760 ;
        RECT 134.420 200.330 135.150 201.680 ;
        RECT 137.640 201.100 137.990 202.930 ;
        RECT 135.870 200.830 137.990 201.100 ;
        RECT 132.550 200.040 133.550 200.050 ;
        RECT 132.110 199.990 132.370 200.010 ;
        RECT 132.540 199.830 133.550 200.040 ;
        RECT 133.690 200.000 135.720 200.330 ;
        RECT 135.880 200.300 136.910 200.830 ;
        RECT 135.895 200.270 136.895 200.300 ;
        RECT 135.895 200.040 136.895 200.060 ;
        RECT 132.540 199.740 133.690 199.830 ;
        RECT 135.870 199.740 136.910 200.040 ;
        RECT 137.070 200.000 137.390 200.330 ;
        RECT 132.540 199.600 136.910 199.740 ;
        RECT 132.540 199.580 135.920 199.600 ;
        RECT 131.490 198.670 133.550 198.940 ;
        RECT 131.490 196.840 131.860 198.670 ;
        RECT 132.110 198.210 132.370 198.240 ;
        RECT 132.110 197.920 132.390 198.210 ;
        RECT 132.550 198.120 133.550 198.670 ;
        RECT 134.420 198.240 135.150 199.580 ;
        RECT 137.640 199.010 137.990 200.830 ;
        RECT 135.870 198.740 137.990 199.010 ;
        RECT 132.550 197.950 133.550 197.960 ;
        RECT 132.110 197.900 132.370 197.920 ;
        RECT 132.540 197.740 133.550 197.950 ;
        RECT 133.690 197.910 135.720 198.240 ;
        RECT 135.880 198.210 136.910 198.740 ;
        RECT 135.895 198.180 136.895 198.210 ;
        RECT 135.895 197.950 136.895 197.970 ;
        RECT 132.540 197.650 133.690 197.740 ;
        RECT 135.870 197.650 136.910 197.950 ;
        RECT 137.070 197.910 137.390 198.240 ;
        RECT 132.540 197.510 136.910 197.650 ;
        RECT 132.540 197.490 135.920 197.510 ;
        RECT 131.490 196.570 133.550 196.840 ;
        RECT 131.490 194.740 131.860 196.570 ;
        RECT 132.110 196.110 132.370 196.140 ;
        RECT 132.110 195.820 132.390 196.110 ;
        RECT 132.550 196.020 133.550 196.570 ;
        RECT 134.420 196.140 135.150 197.490 ;
        RECT 137.640 196.910 137.990 198.740 ;
        RECT 135.870 196.640 137.990 196.910 ;
        RECT 132.550 195.850 133.550 195.860 ;
        RECT 132.110 195.800 132.370 195.820 ;
        RECT 132.540 195.640 133.550 195.850 ;
        RECT 133.690 195.810 135.720 196.140 ;
        RECT 135.880 196.110 136.910 196.640 ;
        RECT 135.895 196.080 136.895 196.110 ;
        RECT 135.895 195.850 136.895 195.870 ;
        RECT 132.540 195.550 133.690 195.640 ;
        RECT 135.870 195.550 136.910 195.850 ;
        RECT 137.070 195.810 137.390 196.140 ;
        RECT 132.540 195.410 136.910 195.550 ;
        RECT 132.540 195.390 135.920 195.410 ;
        RECT 131.490 194.470 133.550 194.740 ;
        RECT 131.490 192.640 131.860 194.470 ;
        RECT 132.110 194.010 132.370 194.040 ;
        RECT 132.110 193.720 132.390 194.010 ;
        RECT 132.550 193.920 133.550 194.470 ;
        RECT 134.420 194.040 135.150 195.390 ;
        RECT 137.640 194.810 137.990 196.640 ;
        RECT 135.870 194.540 137.990 194.810 ;
        RECT 132.550 193.750 133.550 193.760 ;
        RECT 132.110 193.700 132.370 193.720 ;
        RECT 132.540 193.540 133.550 193.750 ;
        RECT 133.690 193.710 135.720 194.040 ;
        RECT 135.880 194.010 136.910 194.540 ;
        RECT 135.895 193.980 136.895 194.010 ;
        RECT 135.895 193.750 136.895 193.770 ;
        RECT 132.540 193.450 133.690 193.540 ;
        RECT 135.870 193.450 136.910 193.750 ;
        RECT 137.070 193.710 137.390 194.040 ;
        RECT 132.540 193.310 136.910 193.450 ;
        RECT 132.540 193.290 135.920 193.310 ;
        RECT 131.490 192.370 133.550 192.640 ;
        RECT 131.490 190.540 131.860 192.370 ;
        RECT 132.110 191.910 132.370 191.940 ;
        RECT 132.110 191.620 132.390 191.910 ;
        RECT 132.550 191.820 133.550 192.370 ;
        RECT 134.420 191.940 135.150 193.290 ;
        RECT 137.640 192.710 137.990 194.540 ;
        RECT 135.870 192.440 137.990 192.710 ;
        RECT 132.550 191.650 133.550 191.660 ;
        RECT 132.110 191.600 132.370 191.620 ;
        RECT 132.540 191.440 133.550 191.650 ;
        RECT 133.690 191.610 135.720 191.940 ;
        RECT 135.880 191.910 136.910 192.440 ;
        RECT 135.895 191.880 136.895 191.910 ;
        RECT 135.895 191.650 136.895 191.670 ;
        RECT 132.540 191.350 133.690 191.440 ;
        RECT 135.870 191.350 136.910 191.650 ;
        RECT 137.070 191.610 137.390 191.940 ;
        RECT 132.540 191.210 136.910 191.350 ;
        RECT 132.540 191.190 135.920 191.210 ;
        RECT 131.490 190.270 133.550 190.540 ;
        RECT 131.490 188.440 131.860 190.270 ;
        RECT 132.110 189.810 132.370 189.840 ;
        RECT 132.110 189.520 132.390 189.810 ;
        RECT 132.550 189.720 133.550 190.270 ;
        RECT 134.420 189.840 135.150 191.190 ;
        RECT 137.640 190.610 137.990 192.440 ;
        RECT 135.870 190.340 137.990 190.610 ;
        RECT 132.550 189.550 133.550 189.560 ;
        RECT 132.110 189.500 132.370 189.520 ;
        RECT 132.540 189.340 133.550 189.550 ;
        RECT 133.690 189.510 135.720 189.840 ;
        RECT 135.880 189.810 136.910 190.340 ;
        RECT 135.895 189.780 136.895 189.810 ;
        RECT 135.895 189.550 136.895 189.570 ;
        RECT 132.540 189.250 133.690 189.340 ;
        RECT 135.870 189.250 136.910 189.550 ;
        RECT 137.070 189.510 137.390 189.840 ;
        RECT 132.540 189.110 136.910 189.250 ;
        RECT 132.540 189.090 135.920 189.110 ;
        RECT 131.490 188.170 133.550 188.440 ;
        RECT 131.490 186.340 131.860 188.170 ;
        RECT 132.110 187.710 132.370 187.740 ;
        RECT 132.110 187.420 132.390 187.710 ;
        RECT 132.550 187.620 133.550 188.170 ;
        RECT 134.420 187.740 135.150 189.090 ;
        RECT 137.640 188.510 137.990 190.340 ;
        RECT 135.870 188.240 137.990 188.510 ;
        RECT 132.550 187.450 133.550 187.460 ;
        RECT 132.110 187.400 132.370 187.420 ;
        RECT 132.540 187.240 133.550 187.450 ;
        RECT 133.690 187.410 135.720 187.740 ;
        RECT 135.880 187.710 136.910 188.240 ;
        RECT 135.895 187.680 136.895 187.710 ;
        RECT 135.895 187.450 136.895 187.470 ;
        RECT 132.540 187.150 133.690 187.240 ;
        RECT 135.870 187.150 136.910 187.450 ;
        RECT 137.070 187.410 137.390 187.740 ;
        RECT 132.540 187.010 136.910 187.150 ;
        RECT 132.540 186.990 135.920 187.010 ;
        RECT 131.490 186.070 133.550 186.340 ;
        RECT 131.490 184.240 131.860 186.070 ;
        RECT 132.110 185.610 132.370 185.640 ;
        RECT 132.110 185.320 132.390 185.610 ;
        RECT 132.550 185.520 133.550 186.070 ;
        RECT 134.420 185.640 135.150 186.990 ;
        RECT 137.640 186.410 137.990 188.240 ;
        RECT 135.870 186.140 137.990 186.410 ;
        RECT 132.550 185.350 133.550 185.360 ;
        RECT 132.110 185.300 132.370 185.320 ;
        RECT 132.540 185.140 133.550 185.350 ;
        RECT 133.690 185.310 135.720 185.640 ;
        RECT 135.880 185.610 136.910 186.140 ;
        RECT 135.895 185.580 136.895 185.610 ;
        RECT 135.895 185.350 136.895 185.370 ;
        RECT 132.540 185.050 133.690 185.140 ;
        RECT 135.870 185.050 136.910 185.350 ;
        RECT 137.070 185.310 137.390 185.640 ;
        RECT 132.540 184.910 136.910 185.050 ;
        RECT 132.540 184.890 135.920 184.910 ;
        RECT 131.490 183.970 133.550 184.240 ;
        RECT 131.490 182.140 131.860 183.970 ;
        RECT 132.110 183.510 132.370 183.540 ;
        RECT 132.110 183.220 132.390 183.510 ;
        RECT 132.550 183.420 133.550 183.970 ;
        RECT 134.420 183.540 135.150 184.890 ;
        RECT 137.640 184.310 137.990 186.140 ;
        RECT 135.870 184.040 137.990 184.310 ;
        RECT 132.550 183.250 133.550 183.260 ;
        RECT 132.110 183.200 132.370 183.220 ;
        RECT 132.540 183.040 133.550 183.250 ;
        RECT 133.690 183.210 135.720 183.540 ;
        RECT 135.880 183.510 136.910 184.040 ;
        RECT 135.895 183.480 136.895 183.510 ;
        RECT 135.895 183.250 136.895 183.270 ;
        RECT 132.540 182.950 133.690 183.040 ;
        RECT 135.870 182.950 136.910 183.250 ;
        RECT 137.070 183.210 137.390 183.540 ;
        RECT 132.540 182.810 136.910 182.950 ;
        RECT 132.540 182.790 135.920 182.810 ;
        RECT 131.490 181.870 133.550 182.140 ;
        RECT 131.490 180.050 131.860 181.870 ;
        RECT 132.110 181.410 132.370 181.440 ;
        RECT 132.110 181.120 132.390 181.410 ;
        RECT 132.550 181.320 133.550 181.870 ;
        RECT 134.420 181.440 135.150 182.790 ;
        RECT 137.640 182.210 137.990 184.040 ;
        RECT 135.870 181.940 137.990 182.210 ;
        RECT 132.550 181.150 133.550 181.160 ;
        RECT 132.110 181.100 132.370 181.120 ;
        RECT 132.540 180.940 133.550 181.150 ;
        RECT 133.690 181.110 135.720 181.440 ;
        RECT 135.880 181.410 136.910 181.940 ;
        RECT 135.895 181.380 136.895 181.410 ;
        RECT 135.895 181.150 136.895 181.170 ;
        RECT 132.540 180.850 133.690 180.940 ;
        RECT 135.870 180.850 136.910 181.150 ;
        RECT 137.070 181.110 137.390 181.440 ;
        RECT 132.540 180.710 136.910 180.850 ;
        RECT 132.540 180.690 135.920 180.710 ;
        RECT 131.490 179.780 133.550 180.050 ;
        RECT 131.490 177.960 131.860 179.780 ;
        RECT 132.110 179.320 132.370 179.350 ;
        RECT 132.110 179.030 132.390 179.320 ;
        RECT 132.550 179.230 133.550 179.780 ;
        RECT 134.420 179.350 135.150 180.690 ;
        RECT 137.640 180.120 137.990 181.940 ;
        RECT 135.870 179.850 137.990 180.120 ;
        RECT 132.550 179.060 133.550 179.070 ;
        RECT 132.110 179.010 132.370 179.030 ;
        RECT 132.540 178.850 133.550 179.060 ;
        RECT 133.690 179.020 135.720 179.350 ;
        RECT 135.880 179.320 136.910 179.850 ;
        RECT 135.895 179.290 136.895 179.320 ;
        RECT 135.895 179.060 136.895 179.080 ;
        RECT 132.540 178.760 133.690 178.850 ;
        RECT 135.870 178.760 136.910 179.060 ;
        RECT 137.070 179.020 137.390 179.350 ;
        RECT 132.540 178.620 136.910 178.760 ;
        RECT 132.540 178.600 135.920 178.620 ;
        RECT 131.490 177.690 133.550 177.960 ;
        RECT 131.490 175.860 131.860 177.690 ;
        RECT 132.110 177.230 132.370 177.260 ;
        RECT 132.110 176.940 132.390 177.230 ;
        RECT 132.550 177.140 133.550 177.690 ;
        RECT 134.420 177.260 135.150 178.600 ;
        RECT 137.640 178.030 137.990 179.850 ;
        RECT 135.870 177.760 137.990 178.030 ;
        RECT 132.550 176.970 133.550 176.980 ;
        RECT 132.110 176.920 132.370 176.940 ;
        RECT 132.540 176.760 133.550 176.970 ;
        RECT 133.690 176.930 135.720 177.260 ;
        RECT 135.880 177.230 136.910 177.760 ;
        RECT 135.895 177.200 136.895 177.230 ;
        RECT 135.895 176.970 136.895 176.990 ;
        RECT 132.540 176.670 133.690 176.760 ;
        RECT 135.870 176.670 136.910 176.970 ;
        RECT 137.070 176.930 137.390 177.260 ;
        RECT 132.540 176.530 136.910 176.670 ;
        RECT 132.540 176.510 135.920 176.530 ;
        RECT 131.490 175.590 133.550 175.860 ;
        RECT 131.490 173.770 131.860 175.590 ;
        RECT 132.110 175.130 132.370 175.160 ;
        RECT 132.110 174.840 132.390 175.130 ;
        RECT 132.550 175.040 133.550 175.590 ;
        RECT 134.420 175.160 135.150 176.510 ;
        RECT 137.640 175.930 137.990 177.760 ;
        RECT 135.870 175.660 137.990 175.930 ;
        RECT 132.550 174.870 133.550 174.880 ;
        RECT 132.110 174.820 132.370 174.840 ;
        RECT 132.540 174.660 133.550 174.870 ;
        RECT 133.690 174.830 135.720 175.160 ;
        RECT 135.880 175.130 136.910 175.660 ;
        RECT 135.895 175.100 136.895 175.130 ;
        RECT 135.895 174.870 136.895 174.890 ;
        RECT 132.540 174.570 133.690 174.660 ;
        RECT 135.870 174.570 136.910 174.870 ;
        RECT 137.070 174.830 137.390 175.160 ;
        RECT 132.540 174.430 136.910 174.570 ;
        RECT 132.540 174.410 135.920 174.430 ;
        RECT 131.490 173.500 133.550 173.770 ;
        RECT 131.490 171.680 131.860 173.500 ;
        RECT 132.110 173.040 132.370 173.070 ;
        RECT 132.110 172.750 132.390 173.040 ;
        RECT 132.550 172.950 133.550 173.500 ;
        RECT 134.420 173.070 135.150 174.410 ;
        RECT 137.640 173.840 137.990 175.660 ;
        RECT 135.870 173.570 137.990 173.840 ;
        RECT 132.550 172.780 133.550 172.790 ;
        RECT 132.110 172.730 132.370 172.750 ;
        RECT 132.540 172.570 133.550 172.780 ;
        RECT 133.690 172.740 135.720 173.070 ;
        RECT 135.880 173.040 136.910 173.570 ;
        RECT 135.895 173.010 136.895 173.040 ;
        RECT 135.895 172.780 136.895 172.800 ;
        RECT 132.540 172.480 133.690 172.570 ;
        RECT 135.870 172.480 136.910 172.780 ;
        RECT 137.070 172.740 137.390 173.070 ;
        RECT 132.540 172.340 136.910 172.480 ;
        RECT 132.540 172.320 135.920 172.340 ;
        RECT 131.490 171.410 133.550 171.680 ;
        RECT 131.490 169.580 131.860 171.410 ;
        RECT 132.110 170.950 132.370 170.980 ;
        RECT 132.110 170.660 132.390 170.950 ;
        RECT 132.550 170.860 133.550 171.410 ;
        RECT 134.420 170.980 135.150 172.320 ;
        RECT 137.640 171.750 137.990 173.570 ;
        RECT 135.870 171.480 137.990 171.750 ;
        RECT 132.550 170.690 133.550 170.700 ;
        RECT 132.110 170.640 132.370 170.660 ;
        RECT 132.540 170.480 133.550 170.690 ;
        RECT 133.690 170.650 135.720 170.980 ;
        RECT 135.880 170.950 136.910 171.480 ;
        RECT 135.895 170.920 136.895 170.950 ;
        RECT 135.895 170.690 136.895 170.710 ;
        RECT 132.540 170.390 133.690 170.480 ;
        RECT 135.870 170.390 136.910 170.690 ;
        RECT 137.070 170.650 137.390 170.980 ;
        RECT 132.540 170.250 136.910 170.390 ;
        RECT 132.540 170.230 135.920 170.250 ;
        RECT 131.490 169.310 133.550 169.580 ;
        RECT 131.490 167.480 131.860 169.310 ;
        RECT 132.110 168.850 132.370 168.880 ;
        RECT 132.110 168.560 132.390 168.850 ;
        RECT 132.550 168.760 133.550 169.310 ;
        RECT 134.420 168.880 135.150 170.230 ;
        RECT 137.640 169.650 137.990 171.480 ;
        RECT 135.870 169.380 137.990 169.650 ;
        RECT 132.550 168.590 133.550 168.600 ;
        RECT 132.110 168.540 132.370 168.560 ;
        RECT 132.540 168.380 133.550 168.590 ;
        RECT 133.690 168.550 135.720 168.880 ;
        RECT 135.880 168.850 136.910 169.380 ;
        RECT 135.895 168.820 136.895 168.850 ;
        RECT 135.895 168.590 136.895 168.610 ;
        RECT 132.540 168.290 133.690 168.380 ;
        RECT 135.870 168.290 136.910 168.590 ;
        RECT 137.070 168.550 137.390 168.880 ;
        RECT 132.540 168.150 136.910 168.290 ;
        RECT 132.540 168.130 135.920 168.150 ;
        RECT 131.490 167.210 133.550 167.480 ;
        RECT 131.490 165.380 131.860 167.210 ;
        RECT 132.110 166.750 132.370 166.780 ;
        RECT 132.110 166.460 132.390 166.750 ;
        RECT 132.550 166.660 133.550 167.210 ;
        RECT 134.420 166.780 135.150 168.130 ;
        RECT 137.640 167.550 137.990 169.380 ;
        RECT 135.870 167.280 137.990 167.550 ;
        RECT 132.550 166.490 133.550 166.500 ;
        RECT 132.110 166.440 132.370 166.460 ;
        RECT 132.540 166.280 133.550 166.490 ;
        RECT 133.690 166.450 135.720 166.780 ;
        RECT 135.880 166.750 136.910 167.280 ;
        RECT 135.895 166.720 136.895 166.750 ;
        RECT 135.895 166.490 136.895 166.510 ;
        RECT 132.540 166.190 133.690 166.280 ;
        RECT 135.870 166.190 136.910 166.490 ;
        RECT 137.070 166.450 137.390 166.780 ;
        RECT 132.540 166.050 136.910 166.190 ;
        RECT 132.540 166.030 135.920 166.050 ;
        RECT 131.490 165.110 133.550 165.380 ;
        RECT 131.490 163.280 131.860 165.110 ;
        RECT 132.110 164.650 132.370 164.680 ;
        RECT 132.110 164.360 132.390 164.650 ;
        RECT 132.550 164.560 133.550 165.110 ;
        RECT 134.420 164.680 135.150 166.030 ;
        RECT 137.640 165.450 137.990 167.280 ;
        RECT 135.870 165.180 137.990 165.450 ;
        RECT 132.550 164.390 133.550 164.400 ;
        RECT 132.110 164.340 132.370 164.360 ;
        RECT 132.540 164.180 133.550 164.390 ;
        RECT 133.690 164.350 135.720 164.680 ;
        RECT 135.880 164.650 136.910 165.180 ;
        RECT 135.895 164.620 136.895 164.650 ;
        RECT 135.895 164.390 136.895 164.410 ;
        RECT 132.540 164.090 133.690 164.180 ;
        RECT 135.870 164.090 136.910 164.390 ;
        RECT 137.070 164.350 137.390 164.680 ;
        RECT 132.540 163.950 136.910 164.090 ;
        RECT 132.540 163.930 135.920 163.950 ;
        RECT 131.490 163.010 133.550 163.280 ;
        RECT 131.490 161.180 131.860 163.010 ;
        RECT 132.110 162.550 132.370 162.580 ;
        RECT 132.110 162.260 132.390 162.550 ;
        RECT 132.550 162.460 133.550 163.010 ;
        RECT 134.420 162.580 135.150 163.930 ;
        RECT 137.640 163.350 137.990 165.180 ;
        RECT 135.870 163.080 137.990 163.350 ;
        RECT 132.550 162.290 133.550 162.300 ;
        RECT 132.110 162.240 132.370 162.260 ;
        RECT 132.540 162.080 133.550 162.290 ;
        RECT 133.690 162.250 135.720 162.580 ;
        RECT 135.880 162.550 136.910 163.080 ;
        RECT 135.895 162.520 136.895 162.550 ;
        RECT 135.895 162.290 136.895 162.310 ;
        RECT 132.540 161.990 133.690 162.080 ;
        RECT 135.870 161.990 136.910 162.290 ;
        RECT 137.070 162.250 137.390 162.580 ;
        RECT 132.540 161.850 136.910 161.990 ;
        RECT 132.540 161.830 135.920 161.850 ;
        RECT 131.490 160.910 133.550 161.180 ;
        RECT 131.490 159.080 131.860 160.910 ;
        RECT 132.110 160.450 132.370 160.480 ;
        RECT 132.110 160.160 132.390 160.450 ;
        RECT 132.550 160.360 133.550 160.910 ;
        RECT 134.420 160.480 135.150 161.830 ;
        RECT 137.640 161.250 137.990 163.080 ;
        RECT 135.870 160.980 137.990 161.250 ;
        RECT 132.550 160.190 133.550 160.200 ;
        RECT 132.110 160.140 132.370 160.160 ;
        RECT 132.540 159.980 133.550 160.190 ;
        RECT 133.690 160.150 135.720 160.480 ;
        RECT 135.880 160.450 136.910 160.980 ;
        RECT 135.895 160.420 136.895 160.450 ;
        RECT 135.895 160.190 136.895 160.210 ;
        RECT 132.540 159.890 133.690 159.980 ;
        RECT 135.870 159.890 136.910 160.190 ;
        RECT 137.070 160.150 137.390 160.480 ;
        RECT 132.540 159.750 136.910 159.890 ;
        RECT 132.540 159.730 135.920 159.750 ;
        RECT 131.490 158.810 133.550 159.080 ;
        RECT 131.490 156.980 131.860 158.810 ;
        RECT 132.110 158.350 132.370 158.380 ;
        RECT 132.110 158.060 132.390 158.350 ;
        RECT 132.550 158.260 133.550 158.810 ;
        RECT 134.420 158.380 135.150 159.730 ;
        RECT 137.640 159.150 137.990 160.980 ;
        RECT 135.870 158.880 137.990 159.150 ;
        RECT 132.550 158.090 133.550 158.100 ;
        RECT 132.110 158.040 132.370 158.060 ;
        RECT 132.540 157.880 133.550 158.090 ;
        RECT 133.690 158.050 135.720 158.380 ;
        RECT 135.880 158.350 136.910 158.880 ;
        RECT 135.895 158.320 136.895 158.350 ;
        RECT 135.895 158.090 136.895 158.110 ;
        RECT 132.540 157.790 133.690 157.880 ;
        RECT 135.870 157.790 136.910 158.090 ;
        RECT 137.070 158.050 137.390 158.380 ;
        RECT 132.540 157.650 136.910 157.790 ;
        RECT 132.540 157.630 135.920 157.650 ;
        RECT 131.490 156.710 133.550 156.980 ;
        RECT 131.490 154.880 131.860 156.710 ;
        RECT 132.110 156.250 132.370 156.280 ;
        RECT 132.110 155.960 132.390 156.250 ;
        RECT 132.550 156.160 133.550 156.710 ;
        RECT 134.420 156.280 135.150 157.630 ;
        RECT 137.640 157.050 137.990 158.880 ;
        RECT 135.870 156.780 137.990 157.050 ;
        RECT 132.550 155.990 133.550 156.000 ;
        RECT 132.110 155.940 132.370 155.960 ;
        RECT 132.540 155.780 133.550 155.990 ;
        RECT 133.690 155.950 135.720 156.280 ;
        RECT 135.880 156.250 136.910 156.780 ;
        RECT 135.895 156.220 136.895 156.250 ;
        RECT 135.895 155.990 136.895 156.010 ;
        RECT 132.540 155.690 133.690 155.780 ;
        RECT 135.870 155.690 136.910 155.990 ;
        RECT 137.070 155.950 137.390 156.280 ;
        RECT 132.540 155.550 136.910 155.690 ;
        RECT 132.540 155.530 135.920 155.550 ;
        RECT 131.490 154.610 133.550 154.880 ;
        RECT 131.490 152.780 131.860 154.610 ;
        RECT 132.110 154.150 132.370 154.180 ;
        RECT 132.110 153.860 132.390 154.150 ;
        RECT 132.550 154.060 133.550 154.610 ;
        RECT 134.420 154.180 135.150 155.530 ;
        RECT 137.640 154.950 137.990 156.780 ;
        RECT 135.870 154.680 137.990 154.950 ;
        RECT 132.550 153.890 133.550 153.900 ;
        RECT 132.110 153.840 132.370 153.860 ;
        RECT 132.540 153.680 133.550 153.890 ;
        RECT 133.690 153.850 135.720 154.180 ;
        RECT 135.880 154.150 136.910 154.680 ;
        RECT 135.895 154.120 136.895 154.150 ;
        RECT 135.895 153.890 136.895 153.910 ;
        RECT 132.540 153.590 133.690 153.680 ;
        RECT 135.870 153.590 136.910 153.890 ;
        RECT 137.070 153.850 137.390 154.180 ;
        RECT 132.540 153.450 136.910 153.590 ;
        RECT 132.540 153.430 135.920 153.450 ;
        RECT 131.490 152.510 133.550 152.780 ;
        RECT 131.490 150.680 131.860 152.510 ;
        RECT 132.110 152.050 132.370 152.080 ;
        RECT 132.110 151.760 132.390 152.050 ;
        RECT 132.550 151.960 133.550 152.510 ;
        RECT 134.420 152.080 135.150 153.430 ;
        RECT 137.640 152.850 137.990 154.680 ;
        RECT 135.870 152.580 137.990 152.850 ;
        RECT 132.550 151.790 133.550 151.800 ;
        RECT 132.110 151.740 132.370 151.760 ;
        RECT 132.540 151.580 133.550 151.790 ;
        RECT 133.690 151.750 135.720 152.080 ;
        RECT 135.880 152.050 136.910 152.580 ;
        RECT 135.895 152.020 136.895 152.050 ;
        RECT 135.895 151.790 136.895 151.810 ;
        RECT 132.540 151.490 133.690 151.580 ;
        RECT 135.870 151.490 136.910 151.790 ;
        RECT 137.070 151.750 137.390 152.080 ;
        RECT 132.540 151.350 136.910 151.490 ;
        RECT 132.540 151.330 135.920 151.350 ;
        RECT 131.490 150.410 133.550 150.680 ;
        RECT 131.490 148.580 131.860 150.410 ;
        RECT 132.110 149.950 132.370 149.980 ;
        RECT 132.110 149.660 132.390 149.950 ;
        RECT 132.550 149.860 133.550 150.410 ;
        RECT 134.420 149.980 135.150 151.330 ;
        RECT 137.640 150.750 137.990 152.580 ;
        RECT 135.870 150.480 137.990 150.750 ;
        RECT 132.550 149.690 133.550 149.700 ;
        RECT 132.110 149.640 132.370 149.660 ;
        RECT 132.540 149.480 133.550 149.690 ;
        RECT 133.690 149.650 135.720 149.980 ;
        RECT 135.880 149.950 136.910 150.480 ;
        RECT 135.895 149.920 136.895 149.950 ;
        RECT 135.895 149.690 136.895 149.710 ;
        RECT 132.540 149.390 133.690 149.480 ;
        RECT 135.870 149.390 136.910 149.690 ;
        RECT 137.070 149.650 137.390 149.980 ;
        RECT 132.540 149.250 136.910 149.390 ;
        RECT 132.540 149.230 135.920 149.250 ;
        RECT 131.490 148.310 133.550 148.580 ;
        RECT 131.490 146.480 131.860 148.310 ;
        RECT 132.110 147.850 132.370 147.880 ;
        RECT 132.110 147.560 132.390 147.850 ;
        RECT 132.550 147.760 133.550 148.310 ;
        RECT 134.420 147.880 135.150 149.230 ;
        RECT 137.640 148.650 137.990 150.480 ;
        RECT 135.870 148.380 137.990 148.650 ;
        RECT 132.550 147.590 133.550 147.600 ;
        RECT 132.110 147.540 132.370 147.560 ;
        RECT 132.540 147.380 133.550 147.590 ;
        RECT 133.690 147.550 135.720 147.880 ;
        RECT 135.880 147.850 136.910 148.380 ;
        RECT 135.895 147.820 136.895 147.850 ;
        RECT 135.895 147.590 136.895 147.610 ;
        RECT 132.540 147.290 133.690 147.380 ;
        RECT 135.870 147.290 136.910 147.590 ;
        RECT 137.070 147.550 137.390 147.880 ;
        RECT 132.540 147.150 136.910 147.290 ;
        RECT 132.540 147.130 135.920 147.150 ;
        RECT 131.490 146.210 133.550 146.480 ;
        RECT 131.490 144.380 131.860 146.210 ;
        RECT 132.110 145.750 132.370 145.780 ;
        RECT 132.110 145.460 132.390 145.750 ;
        RECT 132.550 145.660 133.550 146.210 ;
        RECT 134.420 145.780 135.150 147.130 ;
        RECT 137.640 146.550 137.990 148.380 ;
        RECT 135.870 146.280 137.990 146.550 ;
        RECT 132.550 145.490 133.550 145.500 ;
        RECT 132.110 145.440 132.370 145.460 ;
        RECT 132.540 145.280 133.550 145.490 ;
        RECT 133.690 145.450 135.720 145.780 ;
        RECT 135.880 145.750 136.910 146.280 ;
        RECT 135.895 145.720 136.895 145.750 ;
        RECT 135.895 145.490 136.895 145.510 ;
        RECT 132.540 145.190 133.690 145.280 ;
        RECT 135.870 145.190 136.910 145.490 ;
        RECT 137.070 145.450 137.390 145.780 ;
        RECT 132.540 145.050 136.910 145.190 ;
        RECT 132.540 145.030 135.920 145.050 ;
        RECT 131.490 144.110 133.550 144.380 ;
        RECT 131.490 142.280 131.860 144.110 ;
        RECT 132.110 143.650 132.370 143.680 ;
        RECT 132.110 143.360 132.390 143.650 ;
        RECT 132.550 143.560 133.550 144.110 ;
        RECT 134.420 143.680 135.150 145.030 ;
        RECT 137.640 144.450 137.990 146.280 ;
        RECT 135.870 144.180 137.990 144.450 ;
        RECT 132.550 143.390 133.550 143.400 ;
        RECT 132.110 143.340 132.370 143.360 ;
        RECT 132.540 143.180 133.550 143.390 ;
        RECT 133.690 143.350 135.720 143.680 ;
        RECT 135.880 143.650 136.910 144.180 ;
        RECT 135.895 143.620 136.895 143.650 ;
        RECT 135.895 143.390 136.895 143.410 ;
        RECT 132.540 143.090 133.690 143.180 ;
        RECT 135.870 143.090 136.910 143.390 ;
        RECT 137.070 143.350 137.390 143.680 ;
        RECT 132.540 142.950 136.910 143.090 ;
        RECT 132.540 142.930 135.920 142.950 ;
        RECT 131.490 142.010 133.550 142.280 ;
        RECT 131.490 140.180 131.860 142.010 ;
        RECT 132.110 141.550 132.370 141.580 ;
        RECT 132.110 141.260 132.390 141.550 ;
        RECT 132.550 141.460 133.550 142.010 ;
        RECT 134.420 141.580 135.150 142.930 ;
        RECT 137.640 142.350 137.990 144.180 ;
        RECT 135.870 142.080 137.990 142.350 ;
        RECT 132.550 141.290 133.550 141.300 ;
        RECT 132.110 141.240 132.370 141.260 ;
        RECT 132.540 141.080 133.550 141.290 ;
        RECT 133.690 141.250 135.720 141.580 ;
        RECT 135.880 141.550 136.910 142.080 ;
        RECT 135.895 141.520 136.895 141.550 ;
        RECT 135.895 141.290 136.895 141.310 ;
        RECT 132.540 140.990 133.690 141.080 ;
        RECT 135.870 140.990 136.910 141.290 ;
        RECT 137.070 141.250 137.390 141.580 ;
        RECT 132.540 140.850 136.910 140.990 ;
        RECT 132.540 140.830 135.920 140.850 ;
        RECT 131.490 139.910 133.550 140.180 ;
        RECT 131.490 138.080 131.860 139.910 ;
        RECT 132.110 139.450 132.370 139.480 ;
        RECT 132.110 139.160 132.390 139.450 ;
        RECT 132.550 139.360 133.550 139.910 ;
        RECT 134.420 139.480 135.150 140.830 ;
        RECT 137.640 140.250 137.990 142.080 ;
        RECT 135.870 139.980 137.990 140.250 ;
        RECT 132.550 139.190 133.550 139.200 ;
        RECT 132.110 139.140 132.370 139.160 ;
        RECT 132.540 138.980 133.550 139.190 ;
        RECT 133.690 139.150 135.720 139.480 ;
        RECT 135.880 139.450 136.910 139.980 ;
        RECT 135.895 139.420 136.895 139.450 ;
        RECT 135.895 139.190 136.895 139.210 ;
        RECT 132.540 138.890 133.690 138.980 ;
        RECT 135.870 138.890 136.910 139.190 ;
        RECT 137.070 139.150 137.390 139.480 ;
        RECT 132.540 138.750 136.910 138.890 ;
        RECT 132.540 138.730 135.920 138.750 ;
        RECT 131.490 137.810 133.550 138.080 ;
        RECT 131.490 135.980 131.860 137.810 ;
        RECT 132.110 137.350 132.370 137.380 ;
        RECT 132.110 137.060 132.390 137.350 ;
        RECT 132.550 137.260 133.550 137.810 ;
        RECT 134.420 137.380 135.150 138.730 ;
        RECT 137.640 138.150 137.990 139.980 ;
        RECT 135.870 137.880 137.990 138.150 ;
        RECT 132.550 137.090 133.550 137.100 ;
        RECT 132.110 137.040 132.370 137.060 ;
        RECT 132.540 136.880 133.550 137.090 ;
        RECT 133.690 137.050 135.720 137.380 ;
        RECT 135.880 137.350 136.910 137.880 ;
        RECT 135.895 137.320 136.895 137.350 ;
        RECT 135.895 137.090 136.895 137.110 ;
        RECT 132.540 136.790 133.690 136.880 ;
        RECT 135.870 136.790 136.910 137.090 ;
        RECT 137.070 137.050 137.390 137.380 ;
        RECT 132.540 136.650 136.910 136.790 ;
        RECT 132.540 136.630 135.920 136.650 ;
        RECT 131.490 135.710 133.550 135.980 ;
        RECT 131.490 133.880 131.860 135.710 ;
        RECT 132.110 135.250 132.370 135.280 ;
        RECT 132.110 134.960 132.390 135.250 ;
        RECT 132.550 135.160 133.550 135.710 ;
        RECT 134.420 135.280 135.150 136.630 ;
        RECT 137.640 136.050 137.990 137.880 ;
        RECT 135.870 135.780 137.990 136.050 ;
        RECT 132.550 134.990 133.550 135.000 ;
        RECT 132.110 134.940 132.370 134.960 ;
        RECT 132.540 134.780 133.550 134.990 ;
        RECT 133.690 134.950 135.720 135.280 ;
        RECT 135.880 135.250 136.910 135.780 ;
        RECT 135.895 135.220 136.895 135.250 ;
        RECT 135.895 134.990 136.895 135.010 ;
        RECT 132.540 134.690 133.690 134.780 ;
        RECT 135.870 134.690 136.910 134.990 ;
        RECT 137.070 134.950 137.390 135.280 ;
        RECT 132.540 134.550 136.910 134.690 ;
        RECT 132.540 134.530 135.920 134.550 ;
        RECT 131.490 133.610 133.550 133.880 ;
        RECT 131.490 131.780 131.860 133.610 ;
        RECT 132.110 133.150 132.370 133.180 ;
        RECT 132.110 132.860 132.390 133.150 ;
        RECT 132.550 133.060 133.550 133.610 ;
        RECT 134.420 133.180 135.150 134.530 ;
        RECT 137.640 133.950 137.990 135.780 ;
        RECT 135.870 133.680 137.990 133.950 ;
        RECT 132.550 132.890 133.550 132.900 ;
        RECT 132.110 132.840 132.370 132.860 ;
        RECT 132.540 132.680 133.550 132.890 ;
        RECT 133.690 132.850 135.720 133.180 ;
        RECT 135.880 133.150 136.910 133.680 ;
        RECT 135.895 133.120 136.895 133.150 ;
        RECT 135.895 132.890 136.895 132.910 ;
        RECT 132.540 132.590 133.690 132.680 ;
        RECT 135.870 132.590 136.910 132.890 ;
        RECT 137.070 132.850 137.390 133.180 ;
        RECT 132.540 132.450 136.910 132.590 ;
        RECT 132.540 132.430 135.920 132.450 ;
        RECT 131.490 131.510 133.550 131.780 ;
        RECT 131.490 129.680 131.860 131.510 ;
        RECT 132.110 131.050 132.370 131.080 ;
        RECT 132.110 130.760 132.390 131.050 ;
        RECT 132.550 130.960 133.550 131.510 ;
        RECT 134.420 131.080 135.150 132.430 ;
        RECT 137.640 131.850 137.990 133.680 ;
        RECT 135.870 131.580 137.990 131.850 ;
        RECT 132.550 130.790 133.550 130.800 ;
        RECT 132.110 130.740 132.370 130.760 ;
        RECT 132.540 130.580 133.550 130.790 ;
        RECT 133.690 130.750 135.720 131.080 ;
        RECT 135.880 131.050 136.910 131.580 ;
        RECT 135.895 131.020 136.895 131.050 ;
        RECT 135.895 130.790 136.895 130.810 ;
        RECT 132.540 130.490 133.690 130.580 ;
        RECT 135.870 130.490 136.910 130.790 ;
        RECT 137.070 130.750 137.390 131.080 ;
        RECT 132.540 130.350 136.910 130.490 ;
        RECT 132.540 130.330 135.920 130.350 ;
        RECT 131.490 129.410 133.550 129.680 ;
        RECT 131.490 127.580 131.860 129.410 ;
        RECT 132.110 128.950 132.370 128.980 ;
        RECT 132.110 128.660 132.390 128.950 ;
        RECT 132.550 128.860 133.550 129.410 ;
        RECT 134.420 128.980 135.150 130.330 ;
        RECT 137.640 129.750 137.990 131.580 ;
        RECT 135.870 129.480 137.990 129.750 ;
        RECT 132.550 128.690 133.550 128.700 ;
        RECT 132.110 128.640 132.370 128.660 ;
        RECT 132.540 128.480 133.550 128.690 ;
        RECT 133.690 128.650 135.720 128.980 ;
        RECT 135.880 128.950 136.910 129.480 ;
        RECT 135.895 128.920 136.895 128.950 ;
        RECT 135.895 128.690 136.895 128.710 ;
        RECT 132.540 128.390 133.690 128.480 ;
        RECT 135.870 128.390 136.910 128.690 ;
        RECT 137.070 128.650 137.390 128.980 ;
        RECT 132.540 128.250 136.910 128.390 ;
        RECT 132.540 128.230 135.920 128.250 ;
        RECT 131.490 127.310 133.550 127.580 ;
        RECT 131.490 125.480 131.860 127.310 ;
        RECT 132.110 126.850 132.370 126.880 ;
        RECT 132.110 126.560 132.390 126.850 ;
        RECT 132.550 126.760 133.550 127.310 ;
        RECT 134.420 126.880 135.150 128.230 ;
        RECT 137.640 127.650 137.990 129.480 ;
        RECT 135.870 127.380 137.990 127.650 ;
        RECT 132.550 126.590 133.550 126.600 ;
        RECT 132.110 126.540 132.370 126.560 ;
        RECT 132.540 126.380 133.550 126.590 ;
        RECT 133.690 126.550 135.720 126.880 ;
        RECT 135.880 126.850 136.910 127.380 ;
        RECT 135.895 126.820 136.895 126.850 ;
        RECT 135.895 126.590 136.895 126.610 ;
        RECT 132.540 126.290 133.690 126.380 ;
        RECT 135.870 126.290 136.910 126.590 ;
        RECT 137.070 126.550 137.390 126.880 ;
        RECT 132.540 126.150 136.910 126.290 ;
        RECT 132.540 126.130 135.920 126.150 ;
        RECT 131.490 125.210 133.550 125.480 ;
        RECT 131.490 123.380 131.860 125.210 ;
        RECT 132.110 124.750 132.370 124.780 ;
        RECT 132.110 124.460 132.390 124.750 ;
        RECT 132.550 124.660 133.550 125.210 ;
        RECT 134.420 124.780 135.150 126.130 ;
        RECT 137.640 125.550 137.990 127.380 ;
        RECT 135.870 125.280 137.990 125.550 ;
        RECT 132.550 124.490 133.550 124.500 ;
        RECT 132.110 124.440 132.370 124.460 ;
        RECT 132.540 124.280 133.550 124.490 ;
        RECT 133.690 124.450 135.720 124.780 ;
        RECT 135.880 124.750 136.910 125.280 ;
        RECT 135.895 124.720 136.895 124.750 ;
        RECT 135.895 124.490 136.895 124.510 ;
        RECT 132.540 124.190 133.690 124.280 ;
        RECT 135.870 124.190 136.910 124.490 ;
        RECT 137.070 124.450 137.390 124.780 ;
        RECT 132.540 124.050 136.910 124.190 ;
        RECT 132.540 124.030 135.920 124.050 ;
        RECT 131.490 123.110 133.550 123.380 ;
        RECT 131.490 121.280 131.860 123.110 ;
        RECT 132.110 122.650 132.370 122.680 ;
        RECT 132.110 122.360 132.390 122.650 ;
        RECT 132.550 122.560 133.550 123.110 ;
        RECT 134.420 122.680 135.150 124.030 ;
        RECT 137.640 123.450 137.990 125.280 ;
        RECT 135.870 123.180 137.990 123.450 ;
        RECT 132.550 122.390 133.550 122.400 ;
        RECT 132.110 122.340 132.370 122.360 ;
        RECT 132.540 122.180 133.550 122.390 ;
        RECT 133.690 122.350 135.720 122.680 ;
        RECT 135.880 122.650 136.910 123.180 ;
        RECT 135.895 122.620 136.895 122.650 ;
        RECT 135.895 122.390 136.895 122.410 ;
        RECT 132.540 122.090 133.690 122.180 ;
        RECT 135.870 122.090 136.910 122.390 ;
        RECT 137.070 122.350 137.390 122.680 ;
        RECT 132.540 121.950 136.910 122.090 ;
        RECT 132.540 121.930 135.920 121.950 ;
        RECT 131.490 121.010 133.550 121.280 ;
        RECT 131.490 119.180 131.860 121.010 ;
        RECT 132.110 120.550 132.370 120.580 ;
        RECT 132.110 120.260 132.390 120.550 ;
        RECT 132.550 120.460 133.550 121.010 ;
        RECT 134.420 120.580 135.150 121.930 ;
        RECT 137.640 121.350 137.990 123.180 ;
        RECT 135.870 121.080 137.990 121.350 ;
        RECT 132.550 120.290 133.550 120.300 ;
        RECT 132.110 120.240 132.370 120.260 ;
        RECT 132.540 120.080 133.550 120.290 ;
        RECT 133.690 120.250 135.720 120.580 ;
        RECT 135.880 120.550 136.910 121.080 ;
        RECT 135.895 120.520 136.895 120.550 ;
        RECT 135.895 120.290 136.895 120.310 ;
        RECT 132.540 119.990 133.690 120.080 ;
        RECT 135.870 119.990 136.910 120.290 ;
        RECT 137.070 120.250 137.390 120.580 ;
        RECT 132.540 119.850 136.910 119.990 ;
        RECT 132.540 119.830 135.920 119.850 ;
        RECT 131.490 118.910 133.550 119.180 ;
        RECT 131.490 117.080 131.860 118.910 ;
        RECT 132.110 118.450 132.370 118.480 ;
        RECT 132.110 118.160 132.390 118.450 ;
        RECT 132.550 118.360 133.550 118.910 ;
        RECT 134.420 118.480 135.150 119.830 ;
        RECT 137.640 119.250 137.990 121.080 ;
        RECT 135.870 118.980 137.990 119.250 ;
        RECT 132.550 118.190 133.550 118.200 ;
        RECT 132.110 118.140 132.370 118.160 ;
        RECT 132.540 117.980 133.550 118.190 ;
        RECT 133.690 118.150 135.720 118.480 ;
        RECT 135.880 118.450 136.910 118.980 ;
        RECT 135.895 118.420 136.895 118.450 ;
        RECT 135.895 118.190 136.895 118.210 ;
        RECT 132.540 117.890 133.690 117.980 ;
        RECT 135.870 117.890 136.910 118.190 ;
        RECT 137.070 118.150 137.390 118.480 ;
        RECT 132.540 117.750 136.910 117.890 ;
        RECT 132.540 117.730 135.920 117.750 ;
        RECT 131.490 116.810 133.550 117.080 ;
        RECT 131.490 114.980 131.860 116.810 ;
        RECT 132.110 116.350 132.370 116.380 ;
        RECT 132.110 116.060 132.390 116.350 ;
        RECT 132.550 116.260 133.550 116.810 ;
        RECT 134.420 116.380 135.150 117.730 ;
        RECT 137.640 117.150 137.990 118.980 ;
        RECT 135.870 116.880 137.990 117.150 ;
        RECT 132.550 116.090 133.550 116.100 ;
        RECT 132.110 116.040 132.370 116.060 ;
        RECT 132.540 115.880 133.550 116.090 ;
        RECT 133.690 116.050 135.720 116.380 ;
        RECT 135.880 116.350 136.910 116.880 ;
        RECT 135.895 116.320 136.895 116.350 ;
        RECT 135.895 116.090 136.895 116.110 ;
        RECT 132.540 115.790 133.690 115.880 ;
        RECT 135.870 115.790 136.910 116.090 ;
        RECT 137.070 116.050 137.390 116.380 ;
        RECT 132.540 115.650 136.910 115.790 ;
        RECT 132.540 115.630 135.920 115.650 ;
        RECT 131.490 114.710 133.550 114.980 ;
        RECT 131.490 112.880 131.860 114.710 ;
        RECT 132.110 114.250 132.370 114.280 ;
        RECT 132.110 113.960 132.390 114.250 ;
        RECT 132.550 114.160 133.550 114.710 ;
        RECT 134.420 114.280 135.150 115.630 ;
        RECT 137.640 115.050 137.990 116.880 ;
        RECT 135.870 114.780 137.990 115.050 ;
        RECT 132.550 113.990 133.550 114.000 ;
        RECT 132.110 113.940 132.370 113.960 ;
        RECT 132.540 113.780 133.550 113.990 ;
        RECT 133.690 113.950 135.720 114.280 ;
        RECT 135.880 114.250 136.910 114.780 ;
        RECT 135.895 114.220 136.895 114.250 ;
        RECT 135.895 113.990 136.895 114.010 ;
        RECT 132.540 113.690 133.690 113.780 ;
        RECT 135.870 113.690 136.910 113.990 ;
        RECT 137.070 113.950 137.390 114.280 ;
        RECT 132.540 113.550 136.910 113.690 ;
        RECT 132.540 113.530 135.920 113.550 ;
        RECT 131.490 112.610 133.550 112.880 ;
        RECT 131.490 110.780 131.860 112.610 ;
        RECT 132.110 112.150 132.370 112.180 ;
        RECT 132.110 111.860 132.390 112.150 ;
        RECT 132.550 112.060 133.550 112.610 ;
        RECT 134.420 112.180 135.150 113.530 ;
        RECT 137.640 112.950 137.990 114.780 ;
        RECT 135.870 112.680 137.990 112.950 ;
        RECT 132.550 111.890 133.550 111.900 ;
        RECT 132.110 111.840 132.370 111.860 ;
        RECT 132.540 111.680 133.550 111.890 ;
        RECT 133.690 111.850 135.720 112.180 ;
        RECT 135.880 112.150 136.910 112.680 ;
        RECT 135.895 112.120 136.895 112.150 ;
        RECT 135.895 111.890 136.895 111.910 ;
        RECT 132.540 111.590 133.690 111.680 ;
        RECT 135.870 111.590 136.910 111.890 ;
        RECT 137.070 111.850 137.390 112.180 ;
        RECT 132.540 111.450 136.910 111.590 ;
        RECT 132.540 111.430 135.920 111.450 ;
        RECT 131.490 110.510 133.550 110.780 ;
        RECT 131.490 108.680 131.860 110.510 ;
        RECT 132.110 110.050 132.370 110.080 ;
        RECT 132.110 109.760 132.390 110.050 ;
        RECT 132.550 109.960 133.550 110.510 ;
        RECT 134.420 110.080 135.150 111.430 ;
        RECT 137.640 110.850 137.990 112.680 ;
        RECT 135.870 110.580 137.990 110.850 ;
        RECT 132.550 109.790 133.550 109.800 ;
        RECT 132.110 109.740 132.370 109.760 ;
        RECT 132.540 109.580 133.550 109.790 ;
        RECT 133.690 109.750 135.720 110.080 ;
        RECT 135.880 110.050 136.910 110.580 ;
        RECT 135.895 110.020 136.895 110.050 ;
        RECT 135.895 109.790 136.895 109.810 ;
        RECT 132.540 109.490 133.690 109.580 ;
        RECT 135.870 109.490 136.910 109.790 ;
        RECT 137.070 109.750 137.390 110.080 ;
        RECT 132.540 109.350 136.910 109.490 ;
        RECT 132.540 109.330 135.920 109.350 ;
        RECT 131.490 108.410 133.550 108.680 ;
        RECT 131.490 106.580 131.860 108.410 ;
        RECT 132.110 107.950 132.370 107.980 ;
        RECT 132.110 107.660 132.390 107.950 ;
        RECT 132.550 107.860 133.550 108.410 ;
        RECT 134.420 107.980 135.150 109.330 ;
        RECT 137.640 108.750 137.990 110.580 ;
        RECT 135.870 108.480 137.990 108.750 ;
        RECT 132.550 107.690 133.550 107.700 ;
        RECT 132.110 107.640 132.370 107.660 ;
        RECT 132.540 107.480 133.550 107.690 ;
        RECT 133.690 107.650 135.720 107.980 ;
        RECT 135.880 107.950 136.910 108.480 ;
        RECT 135.895 107.920 136.895 107.950 ;
        RECT 135.895 107.690 136.895 107.710 ;
        RECT 132.540 107.390 133.690 107.480 ;
        RECT 135.870 107.390 136.910 107.690 ;
        RECT 137.070 107.650 137.390 107.980 ;
        RECT 132.540 107.250 136.910 107.390 ;
        RECT 132.540 107.230 135.920 107.250 ;
        RECT 131.490 106.310 133.550 106.580 ;
        RECT 131.490 104.480 131.860 106.310 ;
        RECT 132.110 105.850 132.370 105.880 ;
        RECT 132.110 105.560 132.390 105.850 ;
        RECT 132.550 105.760 133.550 106.310 ;
        RECT 134.420 105.880 135.150 107.230 ;
        RECT 137.640 106.650 137.990 108.480 ;
        RECT 135.870 106.380 137.990 106.650 ;
        RECT 132.550 105.590 133.550 105.600 ;
        RECT 132.110 105.540 132.370 105.560 ;
        RECT 132.540 105.380 133.550 105.590 ;
        RECT 133.690 105.550 135.720 105.880 ;
        RECT 135.880 105.850 136.910 106.380 ;
        RECT 135.895 105.820 136.895 105.850 ;
        RECT 135.895 105.590 136.895 105.610 ;
        RECT 132.540 105.290 133.690 105.380 ;
        RECT 135.870 105.290 136.910 105.590 ;
        RECT 137.070 105.550 137.390 105.880 ;
        RECT 132.540 105.150 136.910 105.290 ;
        RECT 132.540 105.130 135.920 105.150 ;
        RECT 131.490 104.210 133.550 104.480 ;
        RECT 131.490 102.380 131.860 104.210 ;
        RECT 132.110 103.750 132.370 103.780 ;
        RECT 132.110 103.460 132.390 103.750 ;
        RECT 132.550 103.660 133.550 104.210 ;
        RECT 134.420 103.780 135.150 105.130 ;
        RECT 137.640 104.550 137.990 106.380 ;
        RECT 135.870 104.280 137.990 104.550 ;
        RECT 132.550 103.490 133.550 103.500 ;
        RECT 132.110 103.440 132.370 103.460 ;
        RECT 132.540 103.280 133.550 103.490 ;
        RECT 133.690 103.450 135.720 103.780 ;
        RECT 135.880 103.750 136.910 104.280 ;
        RECT 135.895 103.720 136.895 103.750 ;
        RECT 135.895 103.490 136.895 103.510 ;
        RECT 132.540 103.190 133.690 103.280 ;
        RECT 135.870 103.190 136.910 103.490 ;
        RECT 137.070 103.450 137.390 103.780 ;
        RECT 132.540 103.050 136.910 103.190 ;
        RECT 132.540 103.030 135.920 103.050 ;
        RECT 131.490 102.110 133.550 102.380 ;
        RECT 131.490 100.280 131.860 102.110 ;
        RECT 132.110 101.650 132.370 101.680 ;
        RECT 132.110 101.360 132.390 101.650 ;
        RECT 132.550 101.560 133.550 102.110 ;
        RECT 134.420 101.680 135.150 103.030 ;
        RECT 137.640 102.450 137.990 104.280 ;
        RECT 135.870 102.180 137.990 102.450 ;
        RECT 132.550 101.390 133.550 101.400 ;
        RECT 132.110 101.340 132.370 101.360 ;
        RECT 132.540 101.180 133.550 101.390 ;
        RECT 133.690 101.350 135.720 101.680 ;
        RECT 135.880 101.650 136.910 102.180 ;
        RECT 135.895 101.620 136.895 101.650 ;
        RECT 135.895 101.390 136.895 101.410 ;
        RECT 132.540 101.090 133.690 101.180 ;
        RECT 135.870 101.090 136.910 101.390 ;
        RECT 137.070 101.350 137.390 101.680 ;
        RECT 132.540 100.950 136.910 101.090 ;
        RECT 132.540 100.930 135.920 100.950 ;
        RECT 131.490 100.010 133.550 100.280 ;
        RECT 131.490 98.180 131.860 100.010 ;
        RECT 132.110 99.550 132.370 99.580 ;
        RECT 132.110 99.260 132.390 99.550 ;
        RECT 132.550 99.460 133.550 100.010 ;
        RECT 134.420 99.580 135.150 100.930 ;
        RECT 137.640 100.350 137.990 102.180 ;
        RECT 135.870 100.080 137.990 100.350 ;
        RECT 132.550 99.290 133.550 99.300 ;
        RECT 132.110 99.240 132.370 99.260 ;
        RECT 132.540 99.080 133.550 99.290 ;
        RECT 133.690 99.250 135.720 99.580 ;
        RECT 135.880 99.550 136.910 100.080 ;
        RECT 135.895 99.520 136.895 99.550 ;
        RECT 135.895 99.290 136.895 99.310 ;
        RECT 132.540 98.990 133.690 99.080 ;
        RECT 135.870 98.990 136.910 99.290 ;
        RECT 137.070 99.250 137.390 99.580 ;
        RECT 132.540 98.850 136.910 98.990 ;
        RECT 132.540 98.830 135.920 98.850 ;
        RECT 131.490 97.910 133.550 98.180 ;
        RECT 131.490 96.080 131.860 97.910 ;
        RECT 132.110 97.450 132.370 97.480 ;
        RECT 132.110 97.160 132.390 97.450 ;
        RECT 132.550 97.360 133.550 97.910 ;
        RECT 134.420 97.480 135.150 98.830 ;
        RECT 137.640 98.250 137.990 100.080 ;
        RECT 135.870 97.980 137.990 98.250 ;
        RECT 132.550 97.190 133.550 97.200 ;
        RECT 132.110 97.140 132.370 97.160 ;
        RECT 132.540 96.980 133.550 97.190 ;
        RECT 133.690 97.150 135.720 97.480 ;
        RECT 135.880 97.450 136.910 97.980 ;
        RECT 135.895 97.420 136.895 97.450 ;
        RECT 135.895 97.190 136.895 97.210 ;
        RECT 132.540 96.890 133.690 96.980 ;
        RECT 135.870 96.890 136.910 97.190 ;
        RECT 137.070 97.150 137.390 97.480 ;
        RECT 132.540 96.750 136.910 96.890 ;
        RECT 132.540 96.730 135.920 96.750 ;
        RECT 131.490 95.810 133.550 96.080 ;
        RECT 131.490 93.980 131.860 95.810 ;
        RECT 132.110 95.350 132.370 95.380 ;
        RECT 132.110 95.060 132.390 95.350 ;
        RECT 132.550 95.260 133.550 95.810 ;
        RECT 134.420 95.380 135.150 96.730 ;
        RECT 137.640 96.150 137.990 97.980 ;
        RECT 135.870 95.880 137.990 96.150 ;
        RECT 132.550 95.090 133.550 95.100 ;
        RECT 132.110 95.040 132.370 95.060 ;
        RECT 132.540 94.880 133.550 95.090 ;
        RECT 133.690 95.050 135.720 95.380 ;
        RECT 135.880 95.350 136.910 95.880 ;
        RECT 135.895 95.320 136.895 95.350 ;
        RECT 135.895 95.090 136.895 95.110 ;
        RECT 132.540 94.790 133.690 94.880 ;
        RECT 135.870 94.790 136.910 95.090 ;
        RECT 137.070 95.050 137.390 95.380 ;
        RECT 132.540 94.650 136.910 94.790 ;
        RECT 132.540 94.630 135.920 94.650 ;
        RECT 131.490 93.710 133.550 93.980 ;
        RECT 131.490 91.880 131.860 93.710 ;
        RECT 132.110 93.250 132.370 93.280 ;
        RECT 132.110 92.960 132.390 93.250 ;
        RECT 132.550 93.160 133.550 93.710 ;
        RECT 134.420 93.280 135.150 94.630 ;
        RECT 137.640 94.050 137.990 95.880 ;
        RECT 135.870 93.780 137.990 94.050 ;
        RECT 132.550 92.990 133.550 93.000 ;
        RECT 132.110 92.940 132.370 92.960 ;
        RECT 132.540 92.780 133.550 92.990 ;
        RECT 133.690 92.950 135.720 93.280 ;
        RECT 135.880 93.250 136.910 93.780 ;
        RECT 135.895 93.220 136.895 93.250 ;
        RECT 135.895 92.990 136.895 93.010 ;
        RECT 132.540 92.690 133.690 92.780 ;
        RECT 135.870 92.690 136.910 92.990 ;
        RECT 137.070 92.950 137.390 93.280 ;
        RECT 132.540 92.550 136.910 92.690 ;
        RECT 132.540 92.530 135.920 92.550 ;
        RECT 131.490 91.610 133.550 91.880 ;
        RECT 131.490 89.780 131.860 91.610 ;
        RECT 132.110 91.150 132.370 91.180 ;
        RECT 132.110 90.860 132.390 91.150 ;
        RECT 132.550 91.060 133.550 91.610 ;
        RECT 134.420 91.180 135.150 92.530 ;
        RECT 137.640 91.950 137.990 93.780 ;
        RECT 135.870 91.680 137.990 91.950 ;
        RECT 132.550 90.890 133.550 90.900 ;
        RECT 132.110 90.840 132.370 90.860 ;
        RECT 132.540 90.680 133.550 90.890 ;
        RECT 133.690 90.850 135.720 91.180 ;
        RECT 135.880 91.150 136.910 91.680 ;
        RECT 135.895 91.120 136.895 91.150 ;
        RECT 135.895 90.890 136.895 90.910 ;
        RECT 132.540 90.590 133.690 90.680 ;
        RECT 135.870 90.590 136.910 90.890 ;
        RECT 137.070 90.850 137.390 91.180 ;
        RECT 132.540 90.450 136.910 90.590 ;
        RECT 132.540 90.430 135.920 90.450 ;
        RECT 131.490 89.510 133.550 89.780 ;
        RECT 131.490 87.680 131.860 89.510 ;
        RECT 132.110 89.050 132.370 89.080 ;
        RECT 132.110 88.760 132.390 89.050 ;
        RECT 132.550 88.960 133.550 89.510 ;
        RECT 134.420 89.080 135.150 90.430 ;
        RECT 137.640 89.850 137.990 91.680 ;
        RECT 135.870 89.580 137.990 89.850 ;
        RECT 132.550 88.790 133.550 88.800 ;
        RECT 132.110 88.740 132.370 88.760 ;
        RECT 132.540 88.580 133.550 88.790 ;
        RECT 133.690 88.750 135.720 89.080 ;
        RECT 135.880 89.050 136.910 89.580 ;
        RECT 135.895 89.020 136.895 89.050 ;
        RECT 135.895 88.790 136.895 88.810 ;
        RECT 132.540 88.490 133.690 88.580 ;
        RECT 135.870 88.490 136.910 88.790 ;
        RECT 137.070 88.750 137.390 89.080 ;
        RECT 132.540 88.350 136.910 88.490 ;
        RECT 132.540 88.330 135.920 88.350 ;
        RECT 131.490 87.410 133.550 87.680 ;
        RECT 131.490 85.580 131.860 87.410 ;
        RECT 132.110 86.950 132.370 86.980 ;
        RECT 132.110 86.660 132.390 86.950 ;
        RECT 132.550 86.860 133.550 87.410 ;
        RECT 134.420 86.980 135.150 88.330 ;
        RECT 137.640 87.750 137.990 89.580 ;
        RECT 135.870 87.480 137.990 87.750 ;
        RECT 132.550 86.690 133.550 86.700 ;
        RECT 132.110 86.640 132.370 86.660 ;
        RECT 132.540 86.480 133.550 86.690 ;
        RECT 133.690 86.650 135.720 86.980 ;
        RECT 135.880 86.950 136.910 87.480 ;
        RECT 135.895 86.920 136.895 86.950 ;
        RECT 135.895 86.690 136.895 86.710 ;
        RECT 132.540 86.390 133.690 86.480 ;
        RECT 135.870 86.390 136.910 86.690 ;
        RECT 137.070 86.650 137.390 86.980 ;
        RECT 132.540 86.250 136.910 86.390 ;
        RECT 132.540 86.230 135.920 86.250 ;
        RECT 131.490 85.310 133.550 85.580 ;
        RECT 131.490 83.480 131.860 85.310 ;
        RECT 132.110 84.850 132.370 84.880 ;
        RECT 132.110 84.560 132.390 84.850 ;
        RECT 132.550 84.760 133.550 85.310 ;
        RECT 134.420 84.880 135.150 86.230 ;
        RECT 137.640 85.650 137.990 87.480 ;
        RECT 135.870 85.380 137.990 85.650 ;
        RECT 132.550 84.590 133.550 84.600 ;
        RECT 132.110 84.540 132.370 84.560 ;
        RECT 132.540 84.380 133.550 84.590 ;
        RECT 133.690 84.550 135.720 84.880 ;
        RECT 135.880 84.850 136.910 85.380 ;
        RECT 135.895 84.820 136.895 84.850 ;
        RECT 135.895 84.590 136.895 84.610 ;
        RECT 132.540 84.290 133.690 84.380 ;
        RECT 135.870 84.290 136.910 84.590 ;
        RECT 137.070 84.550 137.390 84.880 ;
        RECT 132.540 84.150 136.910 84.290 ;
        RECT 132.540 84.130 135.920 84.150 ;
        RECT 131.490 83.210 133.550 83.480 ;
        RECT 131.490 81.380 131.860 83.210 ;
        RECT 132.110 82.750 132.370 82.780 ;
        RECT 132.110 82.460 132.390 82.750 ;
        RECT 132.550 82.660 133.550 83.210 ;
        RECT 134.420 82.780 135.150 84.130 ;
        RECT 137.640 83.550 137.990 85.380 ;
        RECT 135.870 83.280 137.990 83.550 ;
        RECT 132.550 82.490 133.550 82.500 ;
        RECT 132.110 82.440 132.370 82.460 ;
        RECT 132.540 82.280 133.550 82.490 ;
        RECT 133.690 82.450 135.720 82.780 ;
        RECT 135.880 82.750 136.910 83.280 ;
        RECT 135.895 82.720 136.895 82.750 ;
        RECT 135.895 82.490 136.895 82.510 ;
        RECT 132.540 82.190 133.690 82.280 ;
        RECT 135.870 82.190 136.910 82.490 ;
        RECT 137.070 82.450 137.390 82.780 ;
        RECT 132.540 82.050 136.910 82.190 ;
        RECT 132.540 82.030 135.920 82.050 ;
        RECT 131.490 81.110 133.550 81.380 ;
        RECT 131.490 79.280 131.860 81.110 ;
        RECT 132.110 80.650 132.370 80.680 ;
        RECT 132.110 80.360 132.390 80.650 ;
        RECT 132.550 80.560 133.550 81.110 ;
        RECT 134.420 80.680 135.150 82.030 ;
        RECT 137.640 81.450 137.990 83.280 ;
        RECT 135.870 81.180 137.990 81.450 ;
        RECT 132.550 80.390 133.550 80.400 ;
        RECT 132.110 80.340 132.370 80.360 ;
        RECT 132.540 80.180 133.550 80.390 ;
        RECT 133.690 80.350 135.720 80.680 ;
        RECT 135.880 80.650 136.910 81.180 ;
        RECT 135.895 80.620 136.895 80.650 ;
        RECT 135.895 80.390 136.895 80.410 ;
        RECT 132.540 80.090 133.690 80.180 ;
        RECT 135.870 80.090 136.910 80.390 ;
        RECT 137.070 80.350 137.390 80.680 ;
        RECT 132.540 79.950 136.910 80.090 ;
        RECT 132.540 79.930 135.920 79.950 ;
        RECT 131.490 79.010 133.550 79.280 ;
        RECT 131.490 77.180 131.860 79.010 ;
        RECT 132.110 78.550 132.370 78.580 ;
        RECT 132.110 78.260 132.390 78.550 ;
        RECT 132.550 78.460 133.550 79.010 ;
        RECT 134.420 78.580 135.150 79.930 ;
        RECT 137.640 79.350 137.990 81.180 ;
        RECT 135.870 79.080 137.990 79.350 ;
        RECT 132.550 78.290 133.550 78.300 ;
        RECT 132.110 78.240 132.370 78.260 ;
        RECT 132.540 78.080 133.550 78.290 ;
        RECT 133.690 78.250 135.720 78.580 ;
        RECT 135.880 78.550 136.910 79.080 ;
        RECT 135.895 78.520 136.895 78.550 ;
        RECT 135.895 78.290 136.895 78.310 ;
        RECT 132.540 77.990 133.690 78.080 ;
        RECT 135.870 77.990 136.910 78.290 ;
        RECT 137.070 78.250 137.390 78.580 ;
        RECT 132.540 77.850 136.910 77.990 ;
        RECT 132.540 77.830 135.920 77.850 ;
        RECT 131.490 76.910 133.550 77.180 ;
        RECT 131.490 75.080 131.860 76.910 ;
        RECT 132.110 76.450 132.370 76.480 ;
        RECT 132.110 76.160 132.390 76.450 ;
        RECT 132.550 76.360 133.550 76.910 ;
        RECT 134.420 76.480 135.150 77.830 ;
        RECT 137.640 77.250 137.990 79.080 ;
        RECT 135.870 76.980 137.990 77.250 ;
        RECT 132.550 76.190 133.550 76.200 ;
        RECT 132.110 76.140 132.370 76.160 ;
        RECT 132.540 75.980 133.550 76.190 ;
        RECT 133.690 76.150 135.720 76.480 ;
        RECT 135.880 76.450 136.910 76.980 ;
        RECT 135.895 76.420 136.895 76.450 ;
        RECT 135.895 76.190 136.895 76.210 ;
        RECT 132.540 75.890 133.690 75.980 ;
        RECT 135.870 75.890 136.910 76.190 ;
        RECT 137.070 76.150 137.390 76.480 ;
        RECT 132.540 75.750 136.910 75.890 ;
        RECT 132.540 75.730 135.920 75.750 ;
        RECT 131.490 74.810 133.550 75.080 ;
        RECT 131.490 72.980 131.860 74.810 ;
        RECT 132.110 74.350 132.370 74.380 ;
        RECT 132.110 74.060 132.390 74.350 ;
        RECT 132.550 74.260 133.550 74.810 ;
        RECT 134.420 74.380 135.150 75.730 ;
        RECT 137.640 75.150 137.990 76.980 ;
        RECT 135.870 74.880 137.990 75.150 ;
        RECT 132.550 74.090 133.550 74.100 ;
        RECT 132.110 74.040 132.370 74.060 ;
        RECT 132.540 73.880 133.550 74.090 ;
        RECT 133.690 74.050 135.720 74.380 ;
        RECT 135.880 74.350 136.910 74.880 ;
        RECT 135.895 74.320 136.895 74.350 ;
        RECT 135.895 74.090 136.895 74.110 ;
        RECT 132.540 73.790 133.690 73.880 ;
        RECT 135.870 73.790 136.910 74.090 ;
        RECT 137.070 74.050 137.390 74.380 ;
        RECT 132.540 73.650 136.910 73.790 ;
        RECT 132.540 73.630 135.920 73.650 ;
        RECT 131.490 72.710 133.550 72.980 ;
        RECT 131.490 70.880 131.860 72.710 ;
        RECT 132.110 72.250 132.370 72.280 ;
        RECT 132.110 71.960 132.390 72.250 ;
        RECT 132.550 72.160 133.550 72.710 ;
        RECT 134.420 72.280 135.150 73.630 ;
        RECT 137.640 73.050 137.990 74.880 ;
        RECT 135.870 72.780 137.990 73.050 ;
        RECT 132.550 71.990 133.550 72.000 ;
        RECT 132.110 71.940 132.370 71.960 ;
        RECT 132.540 71.780 133.550 71.990 ;
        RECT 133.690 71.950 135.720 72.280 ;
        RECT 135.880 72.250 136.910 72.780 ;
        RECT 135.895 72.220 136.895 72.250 ;
        RECT 135.895 71.990 136.895 72.010 ;
        RECT 132.540 71.690 133.690 71.780 ;
        RECT 135.870 71.690 136.910 71.990 ;
        RECT 137.070 71.950 137.390 72.280 ;
        RECT 132.540 71.550 136.910 71.690 ;
        RECT 132.540 71.530 135.920 71.550 ;
        RECT 131.490 70.610 133.550 70.880 ;
        RECT 131.490 68.780 131.860 70.610 ;
        RECT 132.110 70.150 132.370 70.180 ;
        RECT 132.110 69.860 132.390 70.150 ;
        RECT 132.550 70.060 133.550 70.610 ;
        RECT 134.420 70.180 135.150 71.530 ;
        RECT 137.640 70.950 137.990 72.780 ;
        RECT 135.870 70.680 137.990 70.950 ;
        RECT 132.550 69.890 133.550 69.900 ;
        RECT 132.110 69.840 132.370 69.860 ;
        RECT 132.540 69.680 133.550 69.890 ;
        RECT 133.690 69.850 135.720 70.180 ;
        RECT 135.880 70.150 136.910 70.680 ;
        RECT 135.895 70.120 136.895 70.150 ;
        RECT 135.895 69.890 136.895 69.910 ;
        RECT 132.540 69.590 133.690 69.680 ;
        RECT 135.870 69.590 136.910 69.890 ;
        RECT 137.070 69.850 137.390 70.180 ;
        RECT 132.540 69.450 136.910 69.590 ;
        RECT 132.540 69.430 135.920 69.450 ;
        RECT 131.490 68.510 133.550 68.780 ;
        RECT 131.490 66.680 131.860 68.510 ;
        RECT 132.110 68.050 132.370 68.080 ;
        RECT 132.110 67.760 132.390 68.050 ;
        RECT 132.550 67.960 133.550 68.510 ;
        RECT 134.420 68.080 135.150 69.430 ;
        RECT 137.640 68.850 137.990 70.680 ;
        RECT 135.870 68.580 137.990 68.850 ;
        RECT 132.550 67.790 133.550 67.800 ;
        RECT 132.110 67.740 132.370 67.760 ;
        RECT 132.540 67.580 133.550 67.790 ;
        RECT 133.690 67.750 135.720 68.080 ;
        RECT 135.880 68.050 136.910 68.580 ;
        RECT 135.895 68.020 136.895 68.050 ;
        RECT 135.895 67.790 136.895 67.810 ;
        RECT 132.540 67.490 133.690 67.580 ;
        RECT 135.870 67.490 136.910 67.790 ;
        RECT 137.070 67.750 137.390 68.080 ;
        RECT 132.540 67.350 136.910 67.490 ;
        RECT 132.540 67.330 135.920 67.350 ;
        RECT 131.490 66.410 133.550 66.680 ;
        RECT 131.490 64.580 131.860 66.410 ;
        RECT 132.110 65.950 132.370 65.980 ;
        RECT 132.110 65.660 132.390 65.950 ;
        RECT 132.550 65.860 133.550 66.410 ;
        RECT 134.420 65.980 135.150 67.330 ;
        RECT 137.640 66.750 137.990 68.580 ;
        RECT 135.870 66.480 137.990 66.750 ;
        RECT 132.550 65.690 133.550 65.700 ;
        RECT 132.110 65.640 132.370 65.660 ;
        RECT 132.540 65.480 133.550 65.690 ;
        RECT 133.690 65.650 135.720 65.980 ;
        RECT 135.880 65.950 136.910 66.480 ;
        RECT 135.895 65.920 136.895 65.950 ;
        RECT 135.895 65.690 136.895 65.710 ;
        RECT 132.540 65.390 133.690 65.480 ;
        RECT 135.870 65.390 136.910 65.690 ;
        RECT 137.070 65.650 137.390 65.980 ;
        RECT 132.540 65.250 136.910 65.390 ;
        RECT 132.540 65.230 135.920 65.250 ;
        RECT 131.490 64.310 133.550 64.580 ;
        RECT 131.490 62.480 131.860 64.310 ;
        RECT 132.110 63.850 132.370 63.880 ;
        RECT 132.110 63.560 132.390 63.850 ;
        RECT 132.550 63.760 133.550 64.310 ;
        RECT 134.420 63.880 135.150 65.230 ;
        RECT 137.640 64.650 137.990 66.480 ;
        RECT 135.870 64.380 137.990 64.650 ;
        RECT 132.550 63.590 133.550 63.600 ;
        RECT 132.110 63.540 132.370 63.560 ;
        RECT 132.540 63.380 133.550 63.590 ;
        RECT 133.690 63.550 135.720 63.880 ;
        RECT 135.880 63.850 136.910 64.380 ;
        RECT 135.895 63.820 136.895 63.850 ;
        RECT 135.895 63.590 136.895 63.610 ;
        RECT 132.540 63.290 133.690 63.380 ;
        RECT 135.870 63.290 136.910 63.590 ;
        RECT 137.070 63.550 137.390 63.880 ;
        RECT 132.540 63.150 136.910 63.290 ;
        RECT 132.540 63.130 135.920 63.150 ;
        RECT 131.490 62.210 133.550 62.480 ;
        RECT 131.490 60.380 131.860 62.210 ;
        RECT 132.110 61.750 132.370 61.780 ;
        RECT 132.110 61.460 132.390 61.750 ;
        RECT 132.550 61.660 133.550 62.210 ;
        RECT 134.420 61.780 135.150 63.130 ;
        RECT 137.640 62.550 137.990 64.380 ;
        RECT 135.870 62.280 137.990 62.550 ;
        RECT 132.550 61.490 133.550 61.500 ;
        RECT 132.110 61.440 132.370 61.460 ;
        RECT 132.540 61.280 133.550 61.490 ;
        RECT 133.690 61.450 135.720 61.780 ;
        RECT 135.880 61.750 136.910 62.280 ;
        RECT 135.895 61.720 136.895 61.750 ;
        RECT 135.895 61.490 136.895 61.510 ;
        RECT 132.540 61.190 133.690 61.280 ;
        RECT 135.870 61.190 136.910 61.490 ;
        RECT 137.070 61.450 137.390 61.780 ;
        RECT 132.540 61.050 136.910 61.190 ;
        RECT 132.540 61.030 135.920 61.050 ;
        RECT 131.490 60.110 133.550 60.380 ;
        RECT 131.490 58.280 131.860 60.110 ;
        RECT 132.110 59.650 132.370 59.680 ;
        RECT 132.110 59.360 132.390 59.650 ;
        RECT 132.550 59.560 133.550 60.110 ;
        RECT 134.420 59.680 135.150 61.030 ;
        RECT 137.640 60.450 137.990 62.280 ;
        RECT 135.870 60.180 137.990 60.450 ;
        RECT 132.550 59.390 133.550 59.400 ;
        RECT 132.110 59.340 132.370 59.360 ;
        RECT 132.540 59.180 133.550 59.390 ;
        RECT 133.690 59.350 135.720 59.680 ;
        RECT 135.880 59.650 136.910 60.180 ;
        RECT 135.895 59.620 136.895 59.650 ;
        RECT 135.895 59.390 136.895 59.410 ;
        RECT 132.540 59.090 133.690 59.180 ;
        RECT 135.870 59.090 136.910 59.390 ;
        RECT 137.070 59.350 137.390 59.680 ;
        RECT 132.540 58.950 136.910 59.090 ;
        RECT 132.540 58.930 135.920 58.950 ;
        RECT 131.490 58.010 133.550 58.280 ;
        RECT 131.490 56.180 131.860 58.010 ;
        RECT 132.110 57.550 132.370 57.580 ;
        RECT 132.110 57.260 132.390 57.550 ;
        RECT 132.550 57.460 133.550 58.010 ;
        RECT 134.420 57.580 135.150 58.930 ;
        RECT 137.640 58.350 137.990 60.180 ;
        RECT 135.870 58.080 137.990 58.350 ;
        RECT 132.550 57.290 133.550 57.300 ;
        RECT 132.110 57.240 132.370 57.260 ;
        RECT 132.540 57.080 133.550 57.290 ;
        RECT 133.690 57.250 135.720 57.580 ;
        RECT 135.880 57.550 136.910 58.080 ;
        RECT 135.895 57.520 136.895 57.550 ;
        RECT 135.895 57.290 136.895 57.310 ;
        RECT 132.540 56.990 133.690 57.080 ;
        RECT 135.870 56.990 136.910 57.290 ;
        RECT 137.070 57.250 137.390 57.580 ;
        RECT 132.540 56.850 136.910 56.990 ;
        RECT 132.540 56.830 135.920 56.850 ;
        RECT 131.490 55.910 133.550 56.180 ;
        RECT 131.490 54.080 131.860 55.910 ;
        RECT 132.110 55.450 132.370 55.480 ;
        RECT 132.110 55.160 132.390 55.450 ;
        RECT 132.550 55.360 133.550 55.910 ;
        RECT 134.420 55.480 135.150 56.830 ;
        RECT 137.640 56.250 137.990 58.080 ;
        RECT 135.870 55.980 137.990 56.250 ;
        RECT 132.550 55.190 133.550 55.200 ;
        RECT 132.110 55.140 132.370 55.160 ;
        RECT 132.540 54.980 133.550 55.190 ;
        RECT 133.690 55.150 135.720 55.480 ;
        RECT 135.880 55.450 136.910 55.980 ;
        RECT 135.895 55.420 136.895 55.450 ;
        RECT 135.895 55.190 136.895 55.210 ;
        RECT 132.540 54.890 133.690 54.980 ;
        RECT 135.870 54.890 136.910 55.190 ;
        RECT 137.070 55.150 137.390 55.480 ;
        RECT 132.540 54.750 136.910 54.890 ;
        RECT 132.540 54.730 135.920 54.750 ;
        RECT 131.490 53.810 133.550 54.080 ;
        RECT 131.490 51.980 131.860 53.810 ;
        RECT 132.110 53.350 132.370 53.380 ;
        RECT 132.110 53.060 132.390 53.350 ;
        RECT 132.550 53.260 133.550 53.810 ;
        RECT 134.420 53.380 135.150 54.730 ;
        RECT 137.640 54.150 137.990 55.980 ;
        RECT 135.870 53.880 137.990 54.150 ;
        RECT 132.550 53.090 133.550 53.100 ;
        RECT 132.110 53.040 132.370 53.060 ;
        RECT 132.540 52.880 133.550 53.090 ;
        RECT 133.690 53.050 135.720 53.380 ;
        RECT 135.880 53.350 136.910 53.880 ;
        RECT 135.895 53.320 136.895 53.350 ;
        RECT 135.895 53.090 136.895 53.110 ;
        RECT 132.540 52.790 133.690 52.880 ;
        RECT 135.870 52.790 136.910 53.090 ;
        RECT 137.070 53.050 137.390 53.380 ;
        RECT 132.540 52.650 136.910 52.790 ;
        RECT 132.540 52.630 135.920 52.650 ;
        RECT 131.490 51.710 133.550 51.980 ;
        RECT 131.490 49.880 131.860 51.710 ;
        RECT 132.110 51.250 132.370 51.280 ;
        RECT 132.110 50.960 132.390 51.250 ;
        RECT 132.550 51.160 133.550 51.710 ;
        RECT 134.420 51.280 135.150 52.630 ;
        RECT 137.640 52.050 137.990 53.880 ;
        RECT 135.870 51.780 137.990 52.050 ;
        RECT 132.550 50.990 133.550 51.000 ;
        RECT 132.110 50.940 132.370 50.960 ;
        RECT 132.540 50.780 133.550 50.990 ;
        RECT 133.690 50.950 135.720 51.280 ;
        RECT 135.880 51.250 136.910 51.780 ;
        RECT 135.895 51.220 136.895 51.250 ;
        RECT 135.895 50.990 136.895 51.010 ;
        RECT 132.540 50.690 133.690 50.780 ;
        RECT 135.870 50.690 136.910 50.990 ;
        RECT 137.070 50.950 137.390 51.280 ;
        RECT 132.540 50.550 136.910 50.690 ;
        RECT 132.540 50.530 135.920 50.550 ;
        RECT 131.490 49.610 133.550 49.880 ;
        RECT 131.490 47.780 131.860 49.610 ;
        RECT 132.110 49.150 132.370 49.180 ;
        RECT 132.110 48.860 132.390 49.150 ;
        RECT 132.550 49.060 133.550 49.610 ;
        RECT 134.420 49.180 135.150 50.530 ;
        RECT 137.640 49.950 137.990 51.780 ;
        RECT 135.870 49.680 137.990 49.950 ;
        RECT 132.550 48.890 133.550 48.900 ;
        RECT 132.110 48.840 132.370 48.860 ;
        RECT 132.540 48.680 133.550 48.890 ;
        RECT 133.690 48.850 135.720 49.180 ;
        RECT 135.880 49.150 136.910 49.680 ;
        RECT 135.895 49.120 136.895 49.150 ;
        RECT 135.895 48.890 136.895 48.910 ;
        RECT 132.540 48.590 133.690 48.680 ;
        RECT 135.870 48.590 136.910 48.890 ;
        RECT 137.070 48.850 137.390 49.180 ;
        RECT 132.540 48.450 136.910 48.590 ;
        RECT 132.540 48.430 135.920 48.450 ;
        RECT 131.490 47.510 133.550 47.780 ;
        RECT 131.490 45.680 131.860 47.510 ;
        RECT 132.110 47.050 132.370 47.080 ;
        RECT 132.110 46.760 132.390 47.050 ;
        RECT 132.550 46.960 133.550 47.510 ;
        RECT 134.420 47.080 135.150 48.430 ;
        RECT 137.640 47.850 137.990 49.680 ;
        RECT 135.870 47.580 137.990 47.850 ;
        RECT 132.550 46.790 133.550 46.800 ;
        RECT 132.110 46.740 132.370 46.760 ;
        RECT 132.540 46.580 133.550 46.790 ;
        RECT 133.690 46.750 135.720 47.080 ;
        RECT 135.880 47.050 136.910 47.580 ;
        RECT 135.895 47.020 136.895 47.050 ;
        RECT 135.895 46.790 136.895 46.810 ;
        RECT 132.540 46.490 133.690 46.580 ;
        RECT 135.870 46.490 136.910 46.790 ;
        RECT 137.070 46.750 137.390 47.080 ;
        RECT 132.540 46.350 136.910 46.490 ;
        RECT 132.540 46.330 135.920 46.350 ;
        RECT 131.490 45.410 133.550 45.680 ;
        RECT 131.490 43.580 131.860 45.410 ;
        RECT 132.110 44.950 132.370 44.980 ;
        RECT 132.110 44.660 132.390 44.950 ;
        RECT 132.550 44.860 133.550 45.410 ;
        RECT 134.420 44.980 135.150 46.330 ;
        RECT 137.640 45.750 137.990 47.580 ;
        RECT 135.870 45.480 137.990 45.750 ;
        RECT 132.550 44.690 133.550 44.700 ;
        RECT 132.110 44.640 132.370 44.660 ;
        RECT 132.540 44.480 133.550 44.690 ;
        RECT 133.690 44.650 135.720 44.980 ;
        RECT 135.880 44.950 136.910 45.480 ;
        RECT 135.895 44.920 136.895 44.950 ;
        RECT 135.895 44.690 136.895 44.710 ;
        RECT 132.540 44.390 133.690 44.480 ;
        RECT 135.870 44.390 136.910 44.690 ;
        RECT 137.070 44.650 137.390 44.980 ;
        RECT 132.540 44.250 136.910 44.390 ;
        RECT 132.540 44.230 135.920 44.250 ;
        RECT 131.490 43.310 133.550 43.580 ;
        RECT 131.490 41.480 131.860 43.310 ;
        RECT 132.110 42.850 132.370 42.880 ;
        RECT 132.110 42.560 132.390 42.850 ;
        RECT 132.550 42.760 133.550 43.310 ;
        RECT 134.420 42.880 135.150 44.230 ;
        RECT 137.640 43.650 137.990 45.480 ;
        RECT 135.870 43.380 137.990 43.650 ;
        RECT 132.550 42.590 133.550 42.600 ;
        RECT 132.110 42.540 132.370 42.560 ;
        RECT 132.540 42.380 133.550 42.590 ;
        RECT 133.690 42.550 135.720 42.880 ;
        RECT 135.880 42.850 136.910 43.380 ;
        RECT 135.895 42.820 136.895 42.850 ;
        RECT 135.895 42.590 136.895 42.610 ;
        RECT 132.540 42.290 133.690 42.380 ;
        RECT 135.870 42.290 136.910 42.590 ;
        RECT 137.070 42.550 137.390 42.880 ;
        RECT 132.540 42.150 136.910 42.290 ;
        RECT 132.540 42.130 135.920 42.150 ;
        RECT 131.490 41.210 133.550 41.480 ;
        RECT 131.490 39.380 131.860 41.210 ;
        RECT 132.110 40.750 132.370 40.780 ;
        RECT 132.110 40.460 132.390 40.750 ;
        RECT 132.550 40.660 133.550 41.210 ;
        RECT 134.420 40.780 135.150 42.130 ;
        RECT 137.640 41.550 137.990 43.380 ;
        RECT 135.870 41.280 137.990 41.550 ;
        RECT 132.550 40.490 133.550 40.500 ;
        RECT 132.110 40.440 132.370 40.460 ;
        RECT 132.540 40.280 133.550 40.490 ;
        RECT 133.690 40.450 135.720 40.780 ;
        RECT 135.880 40.750 136.910 41.280 ;
        RECT 135.895 40.720 136.895 40.750 ;
        RECT 135.895 40.490 136.895 40.510 ;
        RECT 132.540 40.190 133.690 40.280 ;
        RECT 135.870 40.190 136.910 40.490 ;
        RECT 137.070 40.450 137.390 40.780 ;
        RECT 132.540 40.050 136.910 40.190 ;
        RECT 132.540 40.030 135.920 40.050 ;
        RECT 131.490 39.110 133.550 39.380 ;
        RECT 131.490 37.280 131.860 39.110 ;
        RECT 132.110 38.650 132.370 38.680 ;
        RECT 132.110 38.360 132.390 38.650 ;
        RECT 132.550 38.560 133.550 39.110 ;
        RECT 134.420 38.680 135.150 40.030 ;
        RECT 137.640 39.450 137.990 41.280 ;
        RECT 135.870 39.180 137.990 39.450 ;
        RECT 132.550 38.390 133.550 38.400 ;
        RECT 132.110 38.340 132.370 38.360 ;
        RECT 132.540 38.180 133.550 38.390 ;
        RECT 133.690 38.350 135.720 38.680 ;
        RECT 135.880 38.650 136.910 39.180 ;
        RECT 135.895 38.620 136.895 38.650 ;
        RECT 135.895 38.390 136.895 38.410 ;
        RECT 132.540 38.090 133.690 38.180 ;
        RECT 135.870 38.090 136.910 38.390 ;
        RECT 137.070 38.350 137.390 38.680 ;
        RECT 132.540 37.950 136.910 38.090 ;
        RECT 132.540 37.930 135.920 37.950 ;
        RECT 131.490 37.010 133.550 37.280 ;
        RECT 131.490 35.180 131.860 37.010 ;
        RECT 132.110 36.550 132.370 36.580 ;
        RECT 132.110 36.260 132.390 36.550 ;
        RECT 132.550 36.460 133.550 37.010 ;
        RECT 134.420 36.580 135.150 37.930 ;
        RECT 137.640 37.350 137.990 39.180 ;
        RECT 135.870 37.080 137.990 37.350 ;
        RECT 132.550 36.290 133.550 36.300 ;
        RECT 132.110 36.240 132.370 36.260 ;
        RECT 132.540 36.080 133.550 36.290 ;
        RECT 133.690 36.250 135.720 36.580 ;
        RECT 135.880 36.550 136.910 37.080 ;
        RECT 135.895 36.520 136.895 36.550 ;
        RECT 135.895 36.290 136.895 36.310 ;
        RECT 132.540 35.990 133.690 36.080 ;
        RECT 135.870 35.990 136.910 36.290 ;
        RECT 137.070 36.250 137.390 36.580 ;
        RECT 132.540 35.850 136.910 35.990 ;
        RECT 132.540 35.830 135.920 35.850 ;
        RECT 131.490 34.910 133.550 35.180 ;
        RECT 131.490 33.080 131.860 34.910 ;
        RECT 132.110 34.450 132.370 34.480 ;
        RECT 132.110 34.160 132.390 34.450 ;
        RECT 132.550 34.360 133.550 34.910 ;
        RECT 134.420 34.480 135.150 35.830 ;
        RECT 137.640 35.250 137.990 37.080 ;
        RECT 135.870 34.980 137.990 35.250 ;
        RECT 132.550 34.190 133.550 34.200 ;
        RECT 132.110 34.140 132.370 34.160 ;
        RECT 132.540 33.980 133.550 34.190 ;
        RECT 133.690 34.150 135.720 34.480 ;
        RECT 135.880 34.450 136.910 34.980 ;
        RECT 135.895 34.420 136.895 34.450 ;
        RECT 135.895 34.190 136.895 34.210 ;
        RECT 132.540 33.890 133.690 33.980 ;
        RECT 135.870 33.890 136.910 34.190 ;
        RECT 137.070 34.150 137.390 34.480 ;
        RECT 132.540 33.750 136.910 33.890 ;
        RECT 132.540 33.730 135.920 33.750 ;
        RECT 131.490 32.810 133.550 33.080 ;
        RECT 131.490 30.980 131.860 32.810 ;
        RECT 132.110 32.350 132.370 32.380 ;
        RECT 132.110 32.060 132.390 32.350 ;
        RECT 132.550 32.260 133.550 32.810 ;
        RECT 134.420 32.380 135.150 33.730 ;
        RECT 137.640 33.150 137.990 34.980 ;
        RECT 135.870 32.880 137.990 33.150 ;
        RECT 132.550 32.090 133.550 32.100 ;
        RECT 132.110 32.040 132.370 32.060 ;
        RECT 132.540 31.880 133.550 32.090 ;
        RECT 133.690 32.050 135.720 32.380 ;
        RECT 135.880 32.350 136.910 32.880 ;
        RECT 135.895 32.320 136.895 32.350 ;
        RECT 135.895 32.090 136.895 32.110 ;
        RECT 132.540 31.790 133.690 31.880 ;
        RECT 135.870 31.790 136.910 32.090 ;
        RECT 137.070 32.050 137.390 32.380 ;
        RECT 132.540 31.650 136.910 31.790 ;
        RECT 132.540 31.630 135.920 31.650 ;
        RECT 131.490 30.710 133.550 30.980 ;
        RECT 131.490 28.880 131.860 30.710 ;
        RECT 132.110 30.250 132.370 30.280 ;
        RECT 132.110 29.960 132.390 30.250 ;
        RECT 132.550 30.160 133.550 30.710 ;
        RECT 134.420 30.280 135.150 31.630 ;
        RECT 137.640 31.050 137.990 32.880 ;
        RECT 135.870 30.780 137.990 31.050 ;
        RECT 132.550 29.990 133.550 30.000 ;
        RECT 132.110 29.940 132.370 29.960 ;
        RECT 132.540 29.780 133.550 29.990 ;
        RECT 133.690 29.950 135.720 30.280 ;
        RECT 135.880 30.250 136.910 30.780 ;
        RECT 135.895 30.220 136.895 30.250 ;
        RECT 135.895 29.990 136.895 30.010 ;
        RECT 132.540 29.690 133.690 29.780 ;
        RECT 135.870 29.690 136.910 29.990 ;
        RECT 137.070 29.950 137.390 30.280 ;
        RECT 132.540 29.550 136.910 29.690 ;
        RECT 132.540 29.530 135.920 29.550 ;
        RECT 131.490 28.610 133.550 28.880 ;
        RECT 131.490 26.780 131.860 28.610 ;
        RECT 132.110 28.150 132.370 28.180 ;
        RECT 132.110 27.860 132.390 28.150 ;
        RECT 132.550 28.060 133.550 28.610 ;
        RECT 134.420 28.180 135.150 29.530 ;
        RECT 137.640 28.950 137.990 30.780 ;
        RECT 135.870 28.680 137.990 28.950 ;
        RECT 132.550 27.890 133.550 27.900 ;
        RECT 132.110 27.840 132.370 27.860 ;
        RECT 132.540 27.680 133.550 27.890 ;
        RECT 133.690 27.850 135.720 28.180 ;
        RECT 135.880 28.150 136.910 28.680 ;
        RECT 135.895 28.120 136.895 28.150 ;
        RECT 135.895 27.890 136.895 27.910 ;
        RECT 132.540 27.590 133.690 27.680 ;
        RECT 135.870 27.590 136.910 27.890 ;
        RECT 137.070 27.850 137.390 28.180 ;
        RECT 132.540 27.450 136.910 27.590 ;
        RECT 132.540 27.430 135.920 27.450 ;
        RECT 131.490 26.510 133.550 26.780 ;
        RECT 131.490 24.680 131.860 26.510 ;
        RECT 132.110 26.050 132.370 26.080 ;
        RECT 132.110 25.760 132.390 26.050 ;
        RECT 132.550 25.960 133.550 26.510 ;
        RECT 134.420 26.080 135.150 27.430 ;
        RECT 137.640 26.850 137.990 28.680 ;
        RECT 135.870 26.580 137.990 26.850 ;
        RECT 132.550 25.790 133.550 25.800 ;
        RECT 132.110 25.740 132.370 25.760 ;
        RECT 132.540 25.580 133.550 25.790 ;
        RECT 133.690 25.750 135.720 26.080 ;
        RECT 135.880 26.050 136.910 26.580 ;
        RECT 135.895 26.020 136.895 26.050 ;
        RECT 135.895 25.790 136.895 25.810 ;
        RECT 132.540 25.490 133.690 25.580 ;
        RECT 135.870 25.490 136.910 25.790 ;
        RECT 137.070 25.750 137.390 26.080 ;
        RECT 132.540 25.350 136.910 25.490 ;
        RECT 132.540 25.330 135.920 25.350 ;
        RECT 131.490 24.410 133.550 24.680 ;
        RECT 131.490 22.580 131.860 24.410 ;
        RECT 132.110 23.950 132.370 23.980 ;
        RECT 132.110 23.660 132.390 23.950 ;
        RECT 132.550 23.860 133.550 24.410 ;
        RECT 134.420 23.980 135.150 25.330 ;
        RECT 137.640 24.750 137.990 26.580 ;
        RECT 135.870 24.480 137.990 24.750 ;
        RECT 132.550 23.690 133.550 23.700 ;
        RECT 132.110 23.640 132.370 23.660 ;
        RECT 132.540 23.480 133.550 23.690 ;
        RECT 133.690 23.650 135.720 23.980 ;
        RECT 135.880 23.950 136.910 24.480 ;
        RECT 135.895 23.920 136.895 23.950 ;
        RECT 135.895 23.690 136.895 23.710 ;
        RECT 132.540 23.390 133.690 23.480 ;
        RECT 135.870 23.390 136.910 23.690 ;
        RECT 137.070 23.650 137.390 23.980 ;
        RECT 132.540 23.250 136.910 23.390 ;
        RECT 132.540 23.230 135.920 23.250 ;
        RECT 131.490 22.310 133.550 22.580 ;
        RECT 131.490 20.480 131.860 22.310 ;
        RECT 132.110 21.850 132.370 21.880 ;
        RECT 132.110 21.560 132.390 21.850 ;
        RECT 132.550 21.760 133.550 22.310 ;
        RECT 134.420 21.880 135.150 23.230 ;
        RECT 137.640 22.650 137.990 24.480 ;
        RECT 135.870 22.380 137.990 22.650 ;
        RECT 132.550 21.590 133.550 21.600 ;
        RECT 132.110 21.540 132.370 21.560 ;
        RECT 132.540 21.380 133.550 21.590 ;
        RECT 133.690 21.550 135.720 21.880 ;
        RECT 135.880 21.850 136.910 22.380 ;
        RECT 135.895 21.820 136.895 21.850 ;
        RECT 135.895 21.590 136.895 21.610 ;
        RECT 132.540 21.290 133.690 21.380 ;
        RECT 135.870 21.290 136.910 21.590 ;
        RECT 137.070 21.550 137.390 21.880 ;
        RECT 132.540 21.150 136.910 21.290 ;
        RECT 132.540 21.130 135.920 21.150 ;
        RECT 131.490 20.210 133.550 20.480 ;
        RECT 131.490 18.380 131.860 20.210 ;
        RECT 132.110 19.750 132.370 19.780 ;
        RECT 132.110 19.460 132.390 19.750 ;
        RECT 132.550 19.660 133.550 20.210 ;
        RECT 134.420 19.780 135.150 21.130 ;
        RECT 137.640 20.550 137.990 22.380 ;
        RECT 135.870 20.280 137.990 20.550 ;
        RECT 132.550 19.490 133.550 19.500 ;
        RECT 132.110 19.440 132.370 19.460 ;
        RECT 132.540 19.280 133.550 19.490 ;
        RECT 133.690 19.450 135.720 19.780 ;
        RECT 135.880 19.750 136.910 20.280 ;
        RECT 135.895 19.720 136.895 19.750 ;
        RECT 135.895 19.490 136.895 19.510 ;
        RECT 132.540 19.190 133.690 19.280 ;
        RECT 135.870 19.190 136.910 19.490 ;
        RECT 137.070 19.450 137.390 19.780 ;
        RECT 132.540 19.050 136.910 19.190 ;
        RECT 132.540 19.030 135.920 19.050 ;
        RECT 131.490 18.110 133.550 18.380 ;
        RECT 131.490 16.280 131.860 18.110 ;
        RECT 132.110 17.650 132.370 17.680 ;
        RECT 132.110 17.360 132.390 17.650 ;
        RECT 132.550 17.560 133.550 18.110 ;
        RECT 134.420 17.680 135.150 19.030 ;
        RECT 137.640 18.450 137.990 20.280 ;
        RECT 135.870 18.180 137.990 18.450 ;
        RECT 132.550 17.390 133.550 17.400 ;
        RECT 132.110 17.340 132.370 17.360 ;
        RECT 132.540 17.180 133.550 17.390 ;
        RECT 133.690 17.350 135.720 17.680 ;
        RECT 135.880 17.650 136.910 18.180 ;
        RECT 135.895 17.620 136.895 17.650 ;
        RECT 135.895 17.390 136.895 17.410 ;
        RECT 132.540 17.090 133.690 17.180 ;
        RECT 135.870 17.090 136.910 17.390 ;
        RECT 137.070 17.350 137.390 17.680 ;
        RECT 132.540 16.950 136.910 17.090 ;
        RECT 132.540 16.930 135.920 16.950 ;
        RECT 131.490 16.010 133.550 16.280 ;
        RECT 131.490 14.180 131.860 16.010 ;
        RECT 132.110 15.550 132.370 15.580 ;
        RECT 132.110 15.260 132.390 15.550 ;
        RECT 132.550 15.460 133.550 16.010 ;
        RECT 134.420 15.580 135.150 16.930 ;
        RECT 137.640 16.350 137.990 18.180 ;
        RECT 135.870 16.080 137.990 16.350 ;
        RECT 132.550 15.290 133.550 15.300 ;
        RECT 132.110 15.240 132.370 15.260 ;
        RECT 132.540 15.080 133.550 15.290 ;
        RECT 133.690 15.250 135.720 15.580 ;
        RECT 135.880 15.550 136.910 16.080 ;
        RECT 135.895 15.520 136.895 15.550 ;
        RECT 135.895 15.290 136.895 15.310 ;
        RECT 132.540 14.990 133.690 15.080 ;
        RECT 135.870 14.990 136.910 15.290 ;
        RECT 137.070 15.250 137.390 15.580 ;
        RECT 132.540 14.850 136.910 14.990 ;
        RECT 132.540 14.830 135.920 14.850 ;
        RECT 131.490 13.910 133.550 14.180 ;
        RECT 131.490 12.080 131.860 13.910 ;
        RECT 132.110 13.450 132.370 13.480 ;
        RECT 132.110 13.160 132.390 13.450 ;
        RECT 132.550 13.360 133.550 13.910 ;
        RECT 134.420 13.480 135.150 14.830 ;
        RECT 137.640 14.250 137.990 16.080 ;
        RECT 135.870 13.980 137.990 14.250 ;
        RECT 132.550 13.190 133.550 13.200 ;
        RECT 132.110 13.140 132.370 13.160 ;
        RECT 132.540 12.980 133.550 13.190 ;
        RECT 133.690 13.150 135.720 13.480 ;
        RECT 135.880 13.450 136.910 13.980 ;
        RECT 135.895 13.420 136.895 13.450 ;
        RECT 135.895 13.190 136.895 13.210 ;
        RECT 132.540 12.890 133.690 12.980 ;
        RECT 135.870 12.890 136.910 13.190 ;
        RECT 137.070 13.150 137.390 13.480 ;
        RECT 132.540 12.750 136.910 12.890 ;
        RECT 132.540 12.730 135.920 12.750 ;
        RECT 131.490 11.810 133.550 12.080 ;
        RECT 131.490 9.980 131.860 11.810 ;
        RECT 132.110 11.350 132.370 11.380 ;
        RECT 132.110 11.060 132.390 11.350 ;
        RECT 132.550 11.260 133.550 11.810 ;
        RECT 134.420 11.380 135.150 12.730 ;
        RECT 137.640 12.150 137.990 13.980 ;
        RECT 135.870 11.880 137.990 12.150 ;
        RECT 132.550 11.090 133.550 11.100 ;
        RECT 132.110 11.040 132.370 11.060 ;
        RECT 132.540 10.880 133.550 11.090 ;
        RECT 133.690 11.050 135.720 11.380 ;
        RECT 135.880 11.350 136.910 11.880 ;
        RECT 135.895 11.320 136.895 11.350 ;
        RECT 135.895 11.090 136.895 11.110 ;
        RECT 132.540 10.790 133.690 10.880 ;
        RECT 135.870 10.790 136.910 11.090 ;
        RECT 137.070 11.050 137.390 11.380 ;
        RECT 132.540 10.650 136.910 10.790 ;
        RECT 132.540 10.630 135.920 10.650 ;
        RECT 131.490 9.710 133.550 9.980 ;
        RECT 131.490 7.880 131.860 9.710 ;
        RECT 132.110 9.250 132.370 9.280 ;
        RECT 132.110 8.960 132.390 9.250 ;
        RECT 132.550 9.160 133.550 9.710 ;
        RECT 134.420 9.280 135.150 10.630 ;
        RECT 137.640 10.050 137.990 11.880 ;
        RECT 135.870 9.780 137.990 10.050 ;
        RECT 132.550 8.990 133.550 9.000 ;
        RECT 132.110 8.940 132.370 8.960 ;
        RECT 132.540 8.780 133.550 8.990 ;
        RECT 133.690 8.950 135.720 9.280 ;
        RECT 135.880 9.250 136.910 9.780 ;
        RECT 135.895 9.220 136.895 9.250 ;
        RECT 135.895 8.990 136.895 9.010 ;
        RECT 132.540 8.690 133.690 8.780 ;
        RECT 135.870 8.690 136.910 8.990 ;
        RECT 137.070 8.950 137.390 9.280 ;
        RECT 132.540 8.550 136.910 8.690 ;
        RECT 132.540 8.530 135.920 8.550 ;
        RECT 131.490 7.610 133.550 7.880 ;
        RECT 131.490 5.780 131.860 7.610 ;
        RECT 132.110 7.150 132.370 7.180 ;
        RECT 132.110 6.860 132.390 7.150 ;
        RECT 132.550 7.060 133.550 7.610 ;
        RECT 134.420 7.180 135.150 8.530 ;
        RECT 137.640 7.950 137.990 9.780 ;
        RECT 135.870 7.680 137.990 7.950 ;
        RECT 132.550 6.890 133.550 6.900 ;
        RECT 132.110 6.840 132.370 6.860 ;
        RECT 132.540 6.680 133.550 6.890 ;
        RECT 133.690 6.850 135.720 7.180 ;
        RECT 135.880 7.150 136.910 7.680 ;
        RECT 135.895 7.120 136.895 7.150 ;
        RECT 135.895 6.890 136.895 6.910 ;
        RECT 132.540 6.590 133.690 6.680 ;
        RECT 135.870 6.590 136.910 6.890 ;
        RECT 137.070 6.850 137.390 7.180 ;
        RECT 132.540 6.450 136.910 6.590 ;
        RECT 132.540 6.430 135.920 6.450 ;
        RECT 131.490 5.510 133.550 5.780 ;
        RECT 131.490 3.680 131.860 5.510 ;
        RECT 132.110 5.050 132.370 5.080 ;
        RECT 132.110 4.760 132.390 5.050 ;
        RECT 132.550 4.960 133.550 5.510 ;
        RECT 134.420 5.080 135.150 6.430 ;
        RECT 137.640 5.850 137.990 7.680 ;
        RECT 135.870 5.580 137.990 5.850 ;
        RECT 132.550 4.790 133.550 4.800 ;
        RECT 132.110 4.740 132.370 4.760 ;
        RECT 132.540 4.580 133.550 4.790 ;
        RECT 133.690 4.750 135.720 5.080 ;
        RECT 135.880 5.050 136.910 5.580 ;
        RECT 135.895 5.020 136.895 5.050 ;
        RECT 135.895 4.790 136.895 4.810 ;
        RECT 132.540 4.490 133.690 4.580 ;
        RECT 135.870 4.490 136.910 4.790 ;
        RECT 137.070 4.750 137.390 5.080 ;
        RECT 132.540 4.350 136.910 4.490 ;
        RECT 132.540 4.330 135.920 4.350 ;
        RECT 131.490 3.410 133.550 3.680 ;
        RECT 131.490 1.750 131.860 3.410 ;
        RECT 132.110 2.950 132.370 2.980 ;
        RECT 132.110 2.660 132.390 2.950 ;
        RECT 132.550 2.860 133.550 3.410 ;
        RECT 134.420 2.980 135.150 4.330 ;
        RECT 137.640 3.750 137.990 5.580 ;
        RECT 135.870 3.480 137.990 3.750 ;
        RECT 132.550 2.690 133.550 2.700 ;
        RECT 132.110 2.640 132.370 2.660 ;
        RECT 132.540 2.480 133.550 2.690 ;
        RECT 133.690 2.650 135.720 2.980 ;
        RECT 135.880 2.950 136.910 3.480 ;
        RECT 135.895 2.920 136.895 2.950 ;
        RECT 135.895 2.690 136.895 2.710 ;
        RECT 132.540 2.390 133.690 2.480 ;
        RECT 135.870 2.390 136.910 2.690 ;
        RECT 137.070 2.650 137.390 2.980 ;
        RECT 132.540 2.250 136.910 2.390 ;
        RECT 132.540 2.230 135.920 2.250 ;
        RECT 134.420 1.840 135.150 2.230 ;
        RECT 134.410 1.590 135.150 1.840 ;
        RECT 137.640 1.750 137.990 3.480 ;
        RECT 153.540 211.730 153.920 212.010 ;
        RECT 153.540 211.590 153.910 211.730 ;
        RECT 153.540 211.320 155.600 211.590 ;
        RECT 153.540 209.490 153.910 211.320 ;
        RECT 154.160 210.860 154.420 210.890 ;
        RECT 154.160 210.570 154.440 210.860 ;
        RECT 154.600 210.770 155.600 211.320 ;
        RECT 156.470 210.890 157.200 211.760 ;
        RECT 159.690 211.660 160.040 212.420 ;
        RECT 157.920 211.390 160.040 211.660 ;
        RECT 154.600 210.600 155.600 210.610 ;
        RECT 154.160 210.550 154.420 210.570 ;
        RECT 154.590 210.390 155.600 210.600 ;
        RECT 155.740 210.560 157.770 210.890 ;
        RECT 157.930 210.860 158.960 211.390 ;
        RECT 157.945 210.830 158.945 210.860 ;
        RECT 157.945 210.600 158.945 210.620 ;
        RECT 154.590 210.300 155.740 210.390 ;
        RECT 157.920 210.300 158.960 210.600 ;
        RECT 159.120 210.560 159.440 210.890 ;
        RECT 154.590 210.160 158.960 210.300 ;
        RECT 154.590 210.140 157.970 210.160 ;
        RECT 153.540 209.220 155.600 209.490 ;
        RECT 153.540 207.390 153.910 209.220 ;
        RECT 154.160 208.760 154.420 208.790 ;
        RECT 154.160 208.470 154.440 208.760 ;
        RECT 154.600 208.670 155.600 209.220 ;
        RECT 156.470 208.790 157.200 210.140 ;
        RECT 159.690 209.560 160.040 211.390 ;
        RECT 157.920 209.290 160.040 209.560 ;
        RECT 154.600 208.500 155.600 208.510 ;
        RECT 154.160 208.450 154.420 208.470 ;
        RECT 154.590 208.290 155.600 208.500 ;
        RECT 155.740 208.460 157.770 208.790 ;
        RECT 157.930 208.760 158.960 209.290 ;
        RECT 157.945 208.730 158.945 208.760 ;
        RECT 157.945 208.500 158.945 208.520 ;
        RECT 154.590 208.200 155.740 208.290 ;
        RECT 157.920 208.200 158.960 208.500 ;
        RECT 159.120 208.460 159.440 208.790 ;
        RECT 154.590 208.060 158.960 208.200 ;
        RECT 154.590 208.040 157.970 208.060 ;
        RECT 153.540 207.120 155.600 207.390 ;
        RECT 153.540 205.290 153.910 207.120 ;
        RECT 154.160 206.660 154.420 206.690 ;
        RECT 154.160 206.370 154.440 206.660 ;
        RECT 154.600 206.570 155.600 207.120 ;
        RECT 156.470 206.690 157.200 208.040 ;
        RECT 159.690 207.460 160.040 209.290 ;
        RECT 157.920 207.190 160.040 207.460 ;
        RECT 154.600 206.400 155.600 206.410 ;
        RECT 154.160 206.350 154.420 206.370 ;
        RECT 154.590 206.190 155.600 206.400 ;
        RECT 155.740 206.360 157.770 206.690 ;
        RECT 157.930 206.660 158.960 207.190 ;
        RECT 157.945 206.630 158.945 206.660 ;
        RECT 157.945 206.400 158.945 206.420 ;
        RECT 154.590 206.100 155.740 206.190 ;
        RECT 157.920 206.100 158.960 206.400 ;
        RECT 159.120 206.360 159.440 206.690 ;
        RECT 154.590 205.960 158.960 206.100 ;
        RECT 154.590 205.940 157.970 205.960 ;
        RECT 153.540 205.020 155.600 205.290 ;
        RECT 153.540 203.190 153.910 205.020 ;
        RECT 154.160 204.560 154.420 204.590 ;
        RECT 154.160 204.270 154.440 204.560 ;
        RECT 154.600 204.470 155.600 205.020 ;
        RECT 156.470 204.590 157.200 205.940 ;
        RECT 159.690 205.360 160.040 207.190 ;
        RECT 157.920 205.090 160.040 205.360 ;
        RECT 154.600 204.300 155.600 204.310 ;
        RECT 154.160 204.250 154.420 204.270 ;
        RECT 154.590 204.090 155.600 204.300 ;
        RECT 155.740 204.260 157.770 204.590 ;
        RECT 157.930 204.560 158.960 205.090 ;
        RECT 157.945 204.530 158.945 204.560 ;
        RECT 157.945 204.300 158.945 204.320 ;
        RECT 154.590 204.000 155.740 204.090 ;
        RECT 157.920 204.000 158.960 204.300 ;
        RECT 159.120 204.260 159.440 204.590 ;
        RECT 154.590 203.860 158.960 204.000 ;
        RECT 154.590 203.840 157.970 203.860 ;
        RECT 153.540 202.920 155.600 203.190 ;
        RECT 153.540 201.090 153.910 202.920 ;
        RECT 154.160 202.460 154.420 202.490 ;
        RECT 154.160 202.170 154.440 202.460 ;
        RECT 154.600 202.370 155.600 202.920 ;
        RECT 156.470 202.490 157.200 203.840 ;
        RECT 159.690 203.260 160.040 205.090 ;
        RECT 157.920 202.990 160.040 203.260 ;
        RECT 154.600 202.200 155.600 202.210 ;
        RECT 154.160 202.150 154.420 202.170 ;
        RECT 154.590 201.990 155.600 202.200 ;
        RECT 155.740 202.160 157.770 202.490 ;
        RECT 157.930 202.460 158.960 202.990 ;
        RECT 157.945 202.430 158.945 202.460 ;
        RECT 157.945 202.200 158.945 202.220 ;
        RECT 154.590 201.900 155.740 201.990 ;
        RECT 157.920 201.900 158.960 202.200 ;
        RECT 159.120 202.160 159.440 202.490 ;
        RECT 154.590 201.760 158.960 201.900 ;
        RECT 154.590 201.740 157.970 201.760 ;
        RECT 153.540 200.820 155.600 201.090 ;
        RECT 153.540 198.990 153.910 200.820 ;
        RECT 154.160 200.360 154.420 200.390 ;
        RECT 154.160 200.070 154.440 200.360 ;
        RECT 154.600 200.270 155.600 200.820 ;
        RECT 156.470 200.390 157.200 201.740 ;
        RECT 159.690 201.160 160.040 202.990 ;
        RECT 157.920 200.890 160.040 201.160 ;
        RECT 154.600 200.100 155.600 200.110 ;
        RECT 154.160 200.050 154.420 200.070 ;
        RECT 154.590 199.890 155.600 200.100 ;
        RECT 155.740 200.060 157.770 200.390 ;
        RECT 157.930 200.360 158.960 200.890 ;
        RECT 157.945 200.330 158.945 200.360 ;
        RECT 157.945 200.100 158.945 200.120 ;
        RECT 154.590 199.800 155.740 199.890 ;
        RECT 157.920 199.800 158.960 200.100 ;
        RECT 159.120 200.060 159.440 200.390 ;
        RECT 154.590 199.660 158.960 199.800 ;
        RECT 154.590 199.640 157.970 199.660 ;
        RECT 153.540 198.720 155.600 198.990 ;
        RECT 153.540 196.890 153.910 198.720 ;
        RECT 154.160 198.260 154.420 198.290 ;
        RECT 154.160 197.970 154.440 198.260 ;
        RECT 154.600 198.170 155.600 198.720 ;
        RECT 156.470 198.290 157.200 199.640 ;
        RECT 159.690 199.060 160.040 200.890 ;
        RECT 157.920 198.790 160.040 199.060 ;
        RECT 154.600 198.000 155.600 198.010 ;
        RECT 154.160 197.950 154.420 197.970 ;
        RECT 154.590 197.790 155.600 198.000 ;
        RECT 155.740 197.960 157.770 198.290 ;
        RECT 157.930 198.260 158.960 198.790 ;
        RECT 157.945 198.230 158.945 198.260 ;
        RECT 157.945 198.000 158.945 198.020 ;
        RECT 154.590 197.700 155.740 197.790 ;
        RECT 157.920 197.700 158.960 198.000 ;
        RECT 159.120 197.960 159.440 198.290 ;
        RECT 154.590 197.560 158.960 197.700 ;
        RECT 154.590 197.540 157.970 197.560 ;
        RECT 153.540 196.620 155.600 196.890 ;
        RECT 153.540 194.790 153.910 196.620 ;
        RECT 154.160 196.160 154.420 196.190 ;
        RECT 154.160 195.870 154.440 196.160 ;
        RECT 154.600 196.070 155.600 196.620 ;
        RECT 156.470 196.190 157.200 197.540 ;
        RECT 159.690 196.960 160.040 198.790 ;
        RECT 157.920 196.690 160.040 196.960 ;
        RECT 154.600 195.900 155.600 195.910 ;
        RECT 154.160 195.850 154.420 195.870 ;
        RECT 154.590 195.690 155.600 195.900 ;
        RECT 155.740 195.860 157.770 196.190 ;
        RECT 157.930 196.160 158.960 196.690 ;
        RECT 157.945 196.130 158.945 196.160 ;
        RECT 157.945 195.900 158.945 195.920 ;
        RECT 154.590 195.600 155.740 195.690 ;
        RECT 157.920 195.600 158.960 195.900 ;
        RECT 159.120 195.860 159.440 196.190 ;
        RECT 154.590 195.460 158.960 195.600 ;
        RECT 154.590 195.440 157.970 195.460 ;
        RECT 153.540 194.520 155.600 194.790 ;
        RECT 153.540 192.690 153.910 194.520 ;
        RECT 154.160 194.060 154.420 194.090 ;
        RECT 154.160 193.770 154.440 194.060 ;
        RECT 154.600 193.970 155.600 194.520 ;
        RECT 156.470 194.090 157.200 195.440 ;
        RECT 159.690 194.860 160.040 196.690 ;
        RECT 157.920 194.590 160.040 194.860 ;
        RECT 154.600 193.800 155.600 193.810 ;
        RECT 154.160 193.750 154.420 193.770 ;
        RECT 154.590 193.590 155.600 193.800 ;
        RECT 155.740 193.760 157.770 194.090 ;
        RECT 157.930 194.060 158.960 194.590 ;
        RECT 157.945 194.030 158.945 194.060 ;
        RECT 157.945 193.800 158.945 193.820 ;
        RECT 154.590 193.500 155.740 193.590 ;
        RECT 157.920 193.500 158.960 193.800 ;
        RECT 159.120 193.760 159.440 194.090 ;
        RECT 154.590 193.360 158.960 193.500 ;
        RECT 154.590 193.340 157.970 193.360 ;
        RECT 153.540 192.420 155.600 192.690 ;
        RECT 153.540 190.590 153.910 192.420 ;
        RECT 154.160 191.960 154.420 191.990 ;
        RECT 154.160 191.670 154.440 191.960 ;
        RECT 154.600 191.870 155.600 192.420 ;
        RECT 156.470 191.990 157.200 193.340 ;
        RECT 159.690 192.760 160.040 194.590 ;
        RECT 157.920 192.490 160.040 192.760 ;
        RECT 154.600 191.700 155.600 191.710 ;
        RECT 154.160 191.650 154.420 191.670 ;
        RECT 154.590 191.490 155.600 191.700 ;
        RECT 155.740 191.660 157.770 191.990 ;
        RECT 157.930 191.960 158.960 192.490 ;
        RECT 157.945 191.930 158.945 191.960 ;
        RECT 157.945 191.700 158.945 191.720 ;
        RECT 154.590 191.400 155.740 191.490 ;
        RECT 157.920 191.400 158.960 191.700 ;
        RECT 159.120 191.660 159.440 191.990 ;
        RECT 154.590 191.260 158.960 191.400 ;
        RECT 154.590 191.240 157.970 191.260 ;
        RECT 153.540 190.320 155.600 190.590 ;
        RECT 153.540 188.490 153.910 190.320 ;
        RECT 154.160 189.860 154.420 189.890 ;
        RECT 154.160 189.570 154.440 189.860 ;
        RECT 154.600 189.770 155.600 190.320 ;
        RECT 156.470 189.890 157.200 191.240 ;
        RECT 159.690 190.660 160.040 192.490 ;
        RECT 157.920 190.390 160.040 190.660 ;
        RECT 154.600 189.600 155.600 189.610 ;
        RECT 154.160 189.550 154.420 189.570 ;
        RECT 154.590 189.390 155.600 189.600 ;
        RECT 155.740 189.560 157.770 189.890 ;
        RECT 157.930 189.860 158.960 190.390 ;
        RECT 157.945 189.830 158.945 189.860 ;
        RECT 157.945 189.600 158.945 189.620 ;
        RECT 154.590 189.300 155.740 189.390 ;
        RECT 157.920 189.300 158.960 189.600 ;
        RECT 159.120 189.560 159.440 189.890 ;
        RECT 154.590 189.160 158.960 189.300 ;
        RECT 154.590 189.140 157.970 189.160 ;
        RECT 153.540 188.220 155.600 188.490 ;
        RECT 153.540 186.390 153.910 188.220 ;
        RECT 154.160 187.760 154.420 187.790 ;
        RECT 154.160 187.470 154.440 187.760 ;
        RECT 154.600 187.670 155.600 188.220 ;
        RECT 156.470 187.790 157.200 189.140 ;
        RECT 159.690 188.560 160.040 190.390 ;
        RECT 157.920 188.290 160.040 188.560 ;
        RECT 154.600 187.500 155.600 187.510 ;
        RECT 154.160 187.450 154.420 187.470 ;
        RECT 154.590 187.290 155.600 187.500 ;
        RECT 155.740 187.460 157.770 187.790 ;
        RECT 157.930 187.760 158.960 188.290 ;
        RECT 157.945 187.730 158.945 187.760 ;
        RECT 157.945 187.500 158.945 187.520 ;
        RECT 154.590 187.200 155.740 187.290 ;
        RECT 157.920 187.200 158.960 187.500 ;
        RECT 159.120 187.460 159.440 187.790 ;
        RECT 154.590 187.060 158.960 187.200 ;
        RECT 154.590 187.040 157.970 187.060 ;
        RECT 153.540 186.120 155.600 186.390 ;
        RECT 153.540 184.290 153.910 186.120 ;
        RECT 154.160 185.660 154.420 185.690 ;
        RECT 154.160 185.370 154.440 185.660 ;
        RECT 154.600 185.570 155.600 186.120 ;
        RECT 156.470 185.690 157.200 187.040 ;
        RECT 159.690 186.460 160.040 188.290 ;
        RECT 157.920 186.190 160.040 186.460 ;
        RECT 154.600 185.400 155.600 185.410 ;
        RECT 154.160 185.350 154.420 185.370 ;
        RECT 154.590 185.190 155.600 185.400 ;
        RECT 155.740 185.360 157.770 185.690 ;
        RECT 157.930 185.660 158.960 186.190 ;
        RECT 157.945 185.630 158.945 185.660 ;
        RECT 157.945 185.400 158.945 185.420 ;
        RECT 154.590 185.100 155.740 185.190 ;
        RECT 157.920 185.100 158.960 185.400 ;
        RECT 159.120 185.360 159.440 185.690 ;
        RECT 154.590 184.960 158.960 185.100 ;
        RECT 154.590 184.940 157.970 184.960 ;
        RECT 153.540 184.020 155.600 184.290 ;
        RECT 153.540 182.190 153.910 184.020 ;
        RECT 154.160 183.560 154.420 183.590 ;
        RECT 154.160 183.270 154.440 183.560 ;
        RECT 154.600 183.470 155.600 184.020 ;
        RECT 156.470 183.590 157.200 184.940 ;
        RECT 159.690 184.360 160.040 186.190 ;
        RECT 157.920 184.090 160.040 184.360 ;
        RECT 154.600 183.300 155.600 183.310 ;
        RECT 154.160 183.250 154.420 183.270 ;
        RECT 154.590 183.090 155.600 183.300 ;
        RECT 155.740 183.260 157.770 183.590 ;
        RECT 157.930 183.560 158.960 184.090 ;
        RECT 157.945 183.530 158.945 183.560 ;
        RECT 157.945 183.300 158.945 183.320 ;
        RECT 154.590 183.000 155.740 183.090 ;
        RECT 157.920 183.000 158.960 183.300 ;
        RECT 159.120 183.260 159.440 183.590 ;
        RECT 154.590 182.860 158.960 183.000 ;
        RECT 154.590 182.840 157.970 182.860 ;
        RECT 153.540 181.920 155.600 182.190 ;
        RECT 153.540 180.090 153.910 181.920 ;
        RECT 154.160 181.460 154.420 181.490 ;
        RECT 154.160 181.170 154.440 181.460 ;
        RECT 154.600 181.370 155.600 181.920 ;
        RECT 156.470 181.490 157.200 182.840 ;
        RECT 159.690 182.260 160.040 184.090 ;
        RECT 157.920 181.990 160.040 182.260 ;
        RECT 154.600 181.200 155.600 181.210 ;
        RECT 154.160 181.150 154.420 181.170 ;
        RECT 154.590 180.990 155.600 181.200 ;
        RECT 155.740 181.160 157.770 181.490 ;
        RECT 157.930 181.460 158.960 181.990 ;
        RECT 157.945 181.430 158.945 181.460 ;
        RECT 157.945 181.200 158.945 181.220 ;
        RECT 154.590 180.900 155.740 180.990 ;
        RECT 157.920 180.900 158.960 181.200 ;
        RECT 159.120 181.160 159.440 181.490 ;
        RECT 154.590 180.760 158.960 180.900 ;
        RECT 154.590 180.740 157.970 180.760 ;
        RECT 153.540 179.820 155.600 180.090 ;
        RECT 153.540 177.990 153.910 179.820 ;
        RECT 154.160 179.360 154.420 179.390 ;
        RECT 154.160 179.070 154.440 179.360 ;
        RECT 154.600 179.270 155.600 179.820 ;
        RECT 156.470 179.390 157.200 180.740 ;
        RECT 159.690 180.160 160.040 181.990 ;
        RECT 157.920 179.890 160.040 180.160 ;
        RECT 154.600 179.100 155.600 179.110 ;
        RECT 154.160 179.050 154.420 179.070 ;
        RECT 154.590 178.890 155.600 179.100 ;
        RECT 155.740 179.060 157.770 179.390 ;
        RECT 157.930 179.360 158.960 179.890 ;
        RECT 157.945 179.330 158.945 179.360 ;
        RECT 157.945 179.100 158.945 179.120 ;
        RECT 154.590 178.800 155.740 178.890 ;
        RECT 157.920 178.800 158.960 179.100 ;
        RECT 159.120 179.060 159.440 179.390 ;
        RECT 154.590 178.660 158.960 178.800 ;
        RECT 154.590 178.640 157.970 178.660 ;
        RECT 153.540 177.720 155.600 177.990 ;
        RECT 153.540 175.890 153.910 177.720 ;
        RECT 154.160 177.260 154.420 177.290 ;
        RECT 154.160 176.970 154.440 177.260 ;
        RECT 154.600 177.170 155.600 177.720 ;
        RECT 156.470 177.290 157.200 178.640 ;
        RECT 159.690 178.060 160.040 179.890 ;
        RECT 157.920 177.790 160.040 178.060 ;
        RECT 154.600 177.000 155.600 177.010 ;
        RECT 154.160 176.950 154.420 176.970 ;
        RECT 154.590 176.790 155.600 177.000 ;
        RECT 155.740 176.960 157.770 177.290 ;
        RECT 157.930 177.260 158.960 177.790 ;
        RECT 157.945 177.230 158.945 177.260 ;
        RECT 157.945 177.000 158.945 177.020 ;
        RECT 154.590 176.700 155.740 176.790 ;
        RECT 157.920 176.700 158.960 177.000 ;
        RECT 159.120 176.960 159.440 177.290 ;
        RECT 154.590 176.560 158.960 176.700 ;
        RECT 154.590 176.540 157.970 176.560 ;
        RECT 153.540 175.620 155.600 175.890 ;
        RECT 153.540 173.790 153.910 175.620 ;
        RECT 154.160 175.160 154.420 175.190 ;
        RECT 154.160 174.870 154.440 175.160 ;
        RECT 154.600 175.070 155.600 175.620 ;
        RECT 156.470 175.190 157.200 176.540 ;
        RECT 159.690 175.960 160.040 177.790 ;
        RECT 157.920 175.690 160.040 175.960 ;
        RECT 154.600 174.900 155.600 174.910 ;
        RECT 154.160 174.850 154.420 174.870 ;
        RECT 154.590 174.690 155.600 174.900 ;
        RECT 155.740 174.860 157.770 175.190 ;
        RECT 157.930 175.160 158.960 175.690 ;
        RECT 157.945 175.130 158.945 175.160 ;
        RECT 157.945 174.900 158.945 174.920 ;
        RECT 154.590 174.600 155.740 174.690 ;
        RECT 157.920 174.600 158.960 174.900 ;
        RECT 159.120 174.860 159.440 175.190 ;
        RECT 154.590 174.460 158.960 174.600 ;
        RECT 154.590 174.440 157.970 174.460 ;
        RECT 153.540 173.520 155.600 173.790 ;
        RECT 153.540 171.690 153.910 173.520 ;
        RECT 154.160 173.060 154.420 173.090 ;
        RECT 154.160 172.770 154.440 173.060 ;
        RECT 154.600 172.970 155.600 173.520 ;
        RECT 156.470 173.090 157.200 174.440 ;
        RECT 159.690 173.860 160.040 175.690 ;
        RECT 157.920 173.590 160.040 173.860 ;
        RECT 154.600 172.800 155.600 172.810 ;
        RECT 154.160 172.750 154.420 172.770 ;
        RECT 154.590 172.590 155.600 172.800 ;
        RECT 155.740 172.760 157.770 173.090 ;
        RECT 157.930 173.060 158.960 173.590 ;
        RECT 157.945 173.030 158.945 173.060 ;
        RECT 157.945 172.800 158.945 172.820 ;
        RECT 154.590 172.500 155.740 172.590 ;
        RECT 157.920 172.500 158.960 172.800 ;
        RECT 159.120 172.760 159.440 173.090 ;
        RECT 154.590 172.360 158.960 172.500 ;
        RECT 154.590 172.340 157.970 172.360 ;
        RECT 153.540 171.420 155.600 171.690 ;
        RECT 153.540 169.590 153.910 171.420 ;
        RECT 154.160 170.960 154.420 170.990 ;
        RECT 154.160 170.670 154.440 170.960 ;
        RECT 154.600 170.870 155.600 171.420 ;
        RECT 156.470 170.990 157.200 172.340 ;
        RECT 159.690 171.760 160.040 173.590 ;
        RECT 157.920 171.490 160.040 171.760 ;
        RECT 154.600 170.700 155.600 170.710 ;
        RECT 154.160 170.650 154.420 170.670 ;
        RECT 154.590 170.490 155.600 170.700 ;
        RECT 155.740 170.660 157.770 170.990 ;
        RECT 157.930 170.960 158.960 171.490 ;
        RECT 157.945 170.930 158.945 170.960 ;
        RECT 157.945 170.700 158.945 170.720 ;
        RECT 154.590 170.400 155.740 170.490 ;
        RECT 157.920 170.400 158.960 170.700 ;
        RECT 159.120 170.660 159.440 170.990 ;
        RECT 154.590 170.260 158.960 170.400 ;
        RECT 154.590 170.240 157.970 170.260 ;
        RECT 153.540 169.320 155.600 169.590 ;
        RECT 153.540 167.490 153.910 169.320 ;
        RECT 154.160 168.860 154.420 168.890 ;
        RECT 154.160 168.570 154.440 168.860 ;
        RECT 154.600 168.770 155.600 169.320 ;
        RECT 156.470 168.890 157.200 170.240 ;
        RECT 159.690 169.660 160.040 171.490 ;
        RECT 157.920 169.390 160.040 169.660 ;
        RECT 154.600 168.600 155.600 168.610 ;
        RECT 154.160 168.550 154.420 168.570 ;
        RECT 154.590 168.390 155.600 168.600 ;
        RECT 155.740 168.560 157.770 168.890 ;
        RECT 157.930 168.860 158.960 169.390 ;
        RECT 157.945 168.830 158.945 168.860 ;
        RECT 157.945 168.600 158.945 168.620 ;
        RECT 154.590 168.300 155.740 168.390 ;
        RECT 157.920 168.300 158.960 168.600 ;
        RECT 159.120 168.560 159.440 168.890 ;
        RECT 154.590 168.160 158.960 168.300 ;
        RECT 154.590 168.140 157.970 168.160 ;
        RECT 153.540 167.220 155.600 167.490 ;
        RECT 153.540 165.390 153.910 167.220 ;
        RECT 154.160 166.760 154.420 166.790 ;
        RECT 154.160 166.470 154.440 166.760 ;
        RECT 154.600 166.670 155.600 167.220 ;
        RECT 156.470 166.790 157.200 168.140 ;
        RECT 159.690 167.560 160.040 169.390 ;
        RECT 157.920 167.290 160.040 167.560 ;
        RECT 154.600 166.500 155.600 166.510 ;
        RECT 154.160 166.450 154.420 166.470 ;
        RECT 154.590 166.290 155.600 166.500 ;
        RECT 155.740 166.460 157.770 166.790 ;
        RECT 157.930 166.760 158.960 167.290 ;
        RECT 157.945 166.730 158.945 166.760 ;
        RECT 157.945 166.500 158.945 166.520 ;
        RECT 154.590 166.200 155.740 166.290 ;
        RECT 157.920 166.200 158.960 166.500 ;
        RECT 159.120 166.460 159.440 166.790 ;
        RECT 154.590 166.060 158.960 166.200 ;
        RECT 154.590 166.040 157.970 166.060 ;
        RECT 153.540 165.120 155.600 165.390 ;
        RECT 153.540 163.290 153.910 165.120 ;
        RECT 154.160 164.660 154.420 164.690 ;
        RECT 154.160 164.370 154.440 164.660 ;
        RECT 154.600 164.570 155.600 165.120 ;
        RECT 156.470 164.690 157.200 166.040 ;
        RECT 159.690 165.460 160.040 167.290 ;
        RECT 157.920 165.190 160.040 165.460 ;
        RECT 154.600 164.400 155.600 164.410 ;
        RECT 154.160 164.350 154.420 164.370 ;
        RECT 154.590 164.190 155.600 164.400 ;
        RECT 155.740 164.360 157.770 164.690 ;
        RECT 157.930 164.660 158.960 165.190 ;
        RECT 157.945 164.630 158.945 164.660 ;
        RECT 157.945 164.400 158.945 164.420 ;
        RECT 154.590 164.100 155.740 164.190 ;
        RECT 157.920 164.100 158.960 164.400 ;
        RECT 159.120 164.360 159.440 164.690 ;
        RECT 154.590 163.960 158.960 164.100 ;
        RECT 154.590 163.940 157.970 163.960 ;
        RECT 153.540 163.020 155.600 163.290 ;
        RECT 153.540 161.190 153.910 163.020 ;
        RECT 154.160 162.560 154.420 162.590 ;
        RECT 154.160 162.270 154.440 162.560 ;
        RECT 154.600 162.470 155.600 163.020 ;
        RECT 156.470 162.590 157.200 163.940 ;
        RECT 159.690 163.360 160.040 165.190 ;
        RECT 157.920 163.090 160.040 163.360 ;
        RECT 154.600 162.300 155.600 162.310 ;
        RECT 154.160 162.250 154.420 162.270 ;
        RECT 154.590 162.090 155.600 162.300 ;
        RECT 155.740 162.260 157.770 162.590 ;
        RECT 157.930 162.560 158.960 163.090 ;
        RECT 157.945 162.530 158.945 162.560 ;
        RECT 157.945 162.300 158.945 162.320 ;
        RECT 154.590 162.000 155.740 162.090 ;
        RECT 157.920 162.000 158.960 162.300 ;
        RECT 159.120 162.260 159.440 162.590 ;
        RECT 154.590 161.860 158.960 162.000 ;
        RECT 154.590 161.840 157.970 161.860 ;
        RECT 153.540 160.920 155.600 161.190 ;
        RECT 153.540 159.090 153.910 160.920 ;
        RECT 154.160 160.460 154.420 160.490 ;
        RECT 154.160 160.170 154.440 160.460 ;
        RECT 154.600 160.370 155.600 160.920 ;
        RECT 156.470 160.490 157.200 161.840 ;
        RECT 159.690 161.260 160.040 163.090 ;
        RECT 157.920 160.990 160.040 161.260 ;
        RECT 154.600 160.200 155.600 160.210 ;
        RECT 154.160 160.150 154.420 160.170 ;
        RECT 154.590 159.990 155.600 160.200 ;
        RECT 155.740 160.160 157.770 160.490 ;
        RECT 157.930 160.460 158.960 160.990 ;
        RECT 157.945 160.430 158.945 160.460 ;
        RECT 157.945 160.200 158.945 160.220 ;
        RECT 154.590 159.900 155.740 159.990 ;
        RECT 157.920 159.900 158.960 160.200 ;
        RECT 159.120 160.160 159.440 160.490 ;
        RECT 154.590 159.760 158.960 159.900 ;
        RECT 154.590 159.740 157.970 159.760 ;
        RECT 153.540 158.820 155.600 159.090 ;
        RECT 153.540 156.990 153.910 158.820 ;
        RECT 154.160 158.360 154.420 158.390 ;
        RECT 154.160 158.070 154.440 158.360 ;
        RECT 154.600 158.270 155.600 158.820 ;
        RECT 156.470 158.390 157.200 159.740 ;
        RECT 159.690 159.160 160.040 160.990 ;
        RECT 157.920 158.890 160.040 159.160 ;
        RECT 154.600 158.100 155.600 158.110 ;
        RECT 154.160 158.050 154.420 158.070 ;
        RECT 154.590 157.890 155.600 158.100 ;
        RECT 155.740 158.060 157.770 158.390 ;
        RECT 157.930 158.360 158.960 158.890 ;
        RECT 157.945 158.330 158.945 158.360 ;
        RECT 157.945 158.100 158.945 158.120 ;
        RECT 154.590 157.800 155.740 157.890 ;
        RECT 157.920 157.800 158.960 158.100 ;
        RECT 159.120 158.060 159.440 158.390 ;
        RECT 154.590 157.660 158.960 157.800 ;
        RECT 154.590 157.640 157.970 157.660 ;
        RECT 153.540 156.720 155.600 156.990 ;
        RECT 153.540 154.890 153.910 156.720 ;
        RECT 154.160 156.260 154.420 156.290 ;
        RECT 154.160 155.970 154.440 156.260 ;
        RECT 154.600 156.170 155.600 156.720 ;
        RECT 156.470 156.290 157.200 157.640 ;
        RECT 159.690 157.060 160.040 158.890 ;
        RECT 157.920 156.790 160.040 157.060 ;
        RECT 154.600 156.000 155.600 156.010 ;
        RECT 154.160 155.950 154.420 155.970 ;
        RECT 154.590 155.790 155.600 156.000 ;
        RECT 155.740 155.960 157.770 156.290 ;
        RECT 157.930 156.260 158.960 156.790 ;
        RECT 157.945 156.230 158.945 156.260 ;
        RECT 157.945 156.000 158.945 156.020 ;
        RECT 154.590 155.700 155.740 155.790 ;
        RECT 157.920 155.700 158.960 156.000 ;
        RECT 159.120 155.960 159.440 156.290 ;
        RECT 154.590 155.560 158.960 155.700 ;
        RECT 154.590 155.540 157.970 155.560 ;
        RECT 153.540 154.620 155.600 154.890 ;
        RECT 153.540 152.790 153.910 154.620 ;
        RECT 154.160 154.160 154.420 154.190 ;
        RECT 154.160 153.870 154.440 154.160 ;
        RECT 154.600 154.070 155.600 154.620 ;
        RECT 156.470 154.190 157.200 155.540 ;
        RECT 159.690 154.960 160.040 156.790 ;
        RECT 157.920 154.690 160.040 154.960 ;
        RECT 154.600 153.900 155.600 153.910 ;
        RECT 154.160 153.850 154.420 153.870 ;
        RECT 154.590 153.690 155.600 153.900 ;
        RECT 155.740 153.860 157.770 154.190 ;
        RECT 157.930 154.160 158.960 154.690 ;
        RECT 157.945 154.130 158.945 154.160 ;
        RECT 157.945 153.900 158.945 153.920 ;
        RECT 154.590 153.600 155.740 153.690 ;
        RECT 157.920 153.600 158.960 153.900 ;
        RECT 159.120 153.860 159.440 154.190 ;
        RECT 154.590 153.460 158.960 153.600 ;
        RECT 154.590 153.440 157.970 153.460 ;
        RECT 153.540 152.520 155.600 152.790 ;
        RECT 153.540 150.690 153.910 152.520 ;
        RECT 154.160 152.060 154.420 152.090 ;
        RECT 154.160 151.770 154.440 152.060 ;
        RECT 154.600 151.970 155.600 152.520 ;
        RECT 156.470 152.090 157.200 153.440 ;
        RECT 159.690 152.860 160.040 154.690 ;
        RECT 157.920 152.590 160.040 152.860 ;
        RECT 154.600 151.800 155.600 151.810 ;
        RECT 154.160 151.750 154.420 151.770 ;
        RECT 154.590 151.590 155.600 151.800 ;
        RECT 155.740 151.760 157.770 152.090 ;
        RECT 157.930 152.060 158.960 152.590 ;
        RECT 157.945 152.030 158.945 152.060 ;
        RECT 157.945 151.800 158.945 151.820 ;
        RECT 154.590 151.500 155.740 151.590 ;
        RECT 157.920 151.500 158.960 151.800 ;
        RECT 159.120 151.760 159.440 152.090 ;
        RECT 154.590 151.360 158.960 151.500 ;
        RECT 154.590 151.340 157.970 151.360 ;
        RECT 153.540 150.420 155.600 150.690 ;
        RECT 153.540 148.590 153.910 150.420 ;
        RECT 154.160 149.960 154.420 149.990 ;
        RECT 154.160 149.670 154.440 149.960 ;
        RECT 154.600 149.870 155.600 150.420 ;
        RECT 156.470 149.990 157.200 151.340 ;
        RECT 159.690 150.760 160.040 152.590 ;
        RECT 157.920 150.490 160.040 150.760 ;
        RECT 154.600 149.700 155.600 149.710 ;
        RECT 154.160 149.650 154.420 149.670 ;
        RECT 154.590 149.490 155.600 149.700 ;
        RECT 155.740 149.660 157.770 149.990 ;
        RECT 157.930 149.960 158.960 150.490 ;
        RECT 157.945 149.930 158.945 149.960 ;
        RECT 157.945 149.700 158.945 149.720 ;
        RECT 154.590 149.400 155.740 149.490 ;
        RECT 157.920 149.400 158.960 149.700 ;
        RECT 159.120 149.660 159.440 149.990 ;
        RECT 154.590 149.260 158.960 149.400 ;
        RECT 154.590 149.240 157.970 149.260 ;
        RECT 153.540 148.320 155.600 148.590 ;
        RECT 153.540 146.490 153.910 148.320 ;
        RECT 154.160 147.860 154.420 147.890 ;
        RECT 154.160 147.570 154.440 147.860 ;
        RECT 154.600 147.770 155.600 148.320 ;
        RECT 156.470 147.890 157.200 149.240 ;
        RECT 159.690 148.660 160.040 150.490 ;
        RECT 157.920 148.390 160.040 148.660 ;
        RECT 154.600 147.600 155.600 147.610 ;
        RECT 154.160 147.550 154.420 147.570 ;
        RECT 154.590 147.390 155.600 147.600 ;
        RECT 155.740 147.560 157.770 147.890 ;
        RECT 157.930 147.860 158.960 148.390 ;
        RECT 157.945 147.830 158.945 147.860 ;
        RECT 157.945 147.600 158.945 147.620 ;
        RECT 154.590 147.300 155.740 147.390 ;
        RECT 157.920 147.300 158.960 147.600 ;
        RECT 159.120 147.560 159.440 147.890 ;
        RECT 154.590 147.160 158.960 147.300 ;
        RECT 154.590 147.140 157.970 147.160 ;
        RECT 153.540 146.220 155.600 146.490 ;
        RECT 153.540 144.390 153.910 146.220 ;
        RECT 154.160 145.760 154.420 145.790 ;
        RECT 154.160 145.470 154.440 145.760 ;
        RECT 154.600 145.670 155.600 146.220 ;
        RECT 156.470 145.790 157.200 147.140 ;
        RECT 159.690 146.560 160.040 148.390 ;
        RECT 157.920 146.290 160.040 146.560 ;
        RECT 154.600 145.500 155.600 145.510 ;
        RECT 154.160 145.450 154.420 145.470 ;
        RECT 154.590 145.290 155.600 145.500 ;
        RECT 155.740 145.460 157.770 145.790 ;
        RECT 157.930 145.760 158.960 146.290 ;
        RECT 157.945 145.730 158.945 145.760 ;
        RECT 157.945 145.500 158.945 145.520 ;
        RECT 154.590 145.200 155.740 145.290 ;
        RECT 157.920 145.200 158.960 145.500 ;
        RECT 159.120 145.460 159.440 145.790 ;
        RECT 154.590 145.060 158.960 145.200 ;
        RECT 154.590 145.040 157.970 145.060 ;
        RECT 153.540 144.120 155.600 144.390 ;
        RECT 153.540 142.290 153.910 144.120 ;
        RECT 154.160 143.660 154.420 143.690 ;
        RECT 154.160 143.370 154.440 143.660 ;
        RECT 154.600 143.570 155.600 144.120 ;
        RECT 156.470 143.690 157.200 145.040 ;
        RECT 159.690 144.460 160.040 146.290 ;
        RECT 157.920 144.190 160.040 144.460 ;
        RECT 154.600 143.400 155.600 143.410 ;
        RECT 154.160 143.350 154.420 143.370 ;
        RECT 154.590 143.190 155.600 143.400 ;
        RECT 155.740 143.360 157.770 143.690 ;
        RECT 157.930 143.660 158.960 144.190 ;
        RECT 157.945 143.630 158.945 143.660 ;
        RECT 157.945 143.400 158.945 143.420 ;
        RECT 154.590 143.100 155.740 143.190 ;
        RECT 157.920 143.100 158.960 143.400 ;
        RECT 159.120 143.360 159.440 143.690 ;
        RECT 154.590 142.960 158.960 143.100 ;
        RECT 154.590 142.940 157.970 142.960 ;
        RECT 153.540 142.020 155.600 142.290 ;
        RECT 153.540 140.190 153.910 142.020 ;
        RECT 154.160 141.560 154.420 141.590 ;
        RECT 154.160 141.270 154.440 141.560 ;
        RECT 154.600 141.470 155.600 142.020 ;
        RECT 156.470 141.590 157.200 142.940 ;
        RECT 159.690 142.360 160.040 144.190 ;
        RECT 157.920 142.090 160.040 142.360 ;
        RECT 154.600 141.300 155.600 141.310 ;
        RECT 154.160 141.250 154.420 141.270 ;
        RECT 154.590 141.090 155.600 141.300 ;
        RECT 155.740 141.260 157.770 141.590 ;
        RECT 157.930 141.560 158.960 142.090 ;
        RECT 157.945 141.530 158.945 141.560 ;
        RECT 157.945 141.300 158.945 141.320 ;
        RECT 154.590 141.000 155.740 141.090 ;
        RECT 157.920 141.000 158.960 141.300 ;
        RECT 159.120 141.260 159.440 141.590 ;
        RECT 154.590 140.860 158.960 141.000 ;
        RECT 154.590 140.840 157.970 140.860 ;
        RECT 153.540 139.920 155.600 140.190 ;
        RECT 153.540 138.090 153.910 139.920 ;
        RECT 154.160 139.460 154.420 139.490 ;
        RECT 154.160 139.170 154.440 139.460 ;
        RECT 154.600 139.370 155.600 139.920 ;
        RECT 156.470 139.490 157.200 140.840 ;
        RECT 159.690 140.260 160.040 142.090 ;
        RECT 157.920 139.990 160.040 140.260 ;
        RECT 154.600 139.200 155.600 139.210 ;
        RECT 154.160 139.150 154.420 139.170 ;
        RECT 154.590 138.990 155.600 139.200 ;
        RECT 155.740 139.160 157.770 139.490 ;
        RECT 157.930 139.460 158.960 139.990 ;
        RECT 157.945 139.430 158.945 139.460 ;
        RECT 157.945 139.200 158.945 139.220 ;
        RECT 154.590 138.900 155.740 138.990 ;
        RECT 157.920 138.900 158.960 139.200 ;
        RECT 159.120 139.160 159.440 139.490 ;
        RECT 154.590 138.760 158.960 138.900 ;
        RECT 154.590 138.740 157.970 138.760 ;
        RECT 153.540 137.820 155.600 138.090 ;
        RECT 153.540 135.990 153.910 137.820 ;
        RECT 154.160 137.360 154.420 137.390 ;
        RECT 154.160 137.070 154.440 137.360 ;
        RECT 154.600 137.270 155.600 137.820 ;
        RECT 156.470 137.390 157.200 138.740 ;
        RECT 159.690 138.160 160.040 139.990 ;
        RECT 157.920 137.890 160.040 138.160 ;
        RECT 154.600 137.100 155.600 137.110 ;
        RECT 154.160 137.050 154.420 137.070 ;
        RECT 154.590 136.890 155.600 137.100 ;
        RECT 155.740 137.060 157.770 137.390 ;
        RECT 157.930 137.360 158.960 137.890 ;
        RECT 157.945 137.330 158.945 137.360 ;
        RECT 157.945 137.100 158.945 137.120 ;
        RECT 154.590 136.800 155.740 136.890 ;
        RECT 157.920 136.800 158.960 137.100 ;
        RECT 159.120 137.060 159.440 137.390 ;
        RECT 154.590 136.660 158.960 136.800 ;
        RECT 154.590 136.640 157.970 136.660 ;
        RECT 153.540 135.720 155.600 135.990 ;
        RECT 153.540 133.890 153.910 135.720 ;
        RECT 154.160 135.260 154.420 135.290 ;
        RECT 154.160 134.970 154.440 135.260 ;
        RECT 154.600 135.170 155.600 135.720 ;
        RECT 156.470 135.290 157.200 136.640 ;
        RECT 159.690 136.060 160.040 137.890 ;
        RECT 157.920 135.790 160.040 136.060 ;
        RECT 154.600 135.000 155.600 135.010 ;
        RECT 154.160 134.950 154.420 134.970 ;
        RECT 154.590 134.790 155.600 135.000 ;
        RECT 155.740 134.960 157.770 135.290 ;
        RECT 157.930 135.260 158.960 135.790 ;
        RECT 157.945 135.230 158.945 135.260 ;
        RECT 157.945 135.000 158.945 135.020 ;
        RECT 154.590 134.700 155.740 134.790 ;
        RECT 157.920 134.700 158.960 135.000 ;
        RECT 159.120 134.960 159.440 135.290 ;
        RECT 154.590 134.560 158.960 134.700 ;
        RECT 154.590 134.540 157.970 134.560 ;
        RECT 153.540 133.620 155.600 133.890 ;
        RECT 153.540 131.790 153.910 133.620 ;
        RECT 154.160 133.160 154.420 133.190 ;
        RECT 154.160 132.870 154.440 133.160 ;
        RECT 154.600 133.070 155.600 133.620 ;
        RECT 156.470 133.190 157.200 134.540 ;
        RECT 159.690 133.960 160.040 135.790 ;
        RECT 157.920 133.690 160.040 133.960 ;
        RECT 154.600 132.900 155.600 132.910 ;
        RECT 154.160 132.850 154.420 132.870 ;
        RECT 154.590 132.690 155.600 132.900 ;
        RECT 155.740 132.860 157.770 133.190 ;
        RECT 157.930 133.160 158.960 133.690 ;
        RECT 157.945 133.130 158.945 133.160 ;
        RECT 157.945 132.900 158.945 132.920 ;
        RECT 154.590 132.600 155.740 132.690 ;
        RECT 157.920 132.600 158.960 132.900 ;
        RECT 159.120 132.860 159.440 133.190 ;
        RECT 154.590 132.460 158.960 132.600 ;
        RECT 154.590 132.440 157.970 132.460 ;
        RECT 153.540 131.520 155.600 131.790 ;
        RECT 153.540 129.690 153.910 131.520 ;
        RECT 154.160 131.060 154.420 131.090 ;
        RECT 154.160 130.770 154.440 131.060 ;
        RECT 154.600 130.970 155.600 131.520 ;
        RECT 156.470 131.090 157.200 132.440 ;
        RECT 159.690 131.860 160.040 133.690 ;
        RECT 157.920 131.590 160.040 131.860 ;
        RECT 154.600 130.800 155.600 130.810 ;
        RECT 154.160 130.750 154.420 130.770 ;
        RECT 154.590 130.590 155.600 130.800 ;
        RECT 155.740 130.760 157.770 131.090 ;
        RECT 157.930 131.060 158.960 131.590 ;
        RECT 157.945 131.030 158.945 131.060 ;
        RECT 157.945 130.800 158.945 130.820 ;
        RECT 154.590 130.500 155.740 130.590 ;
        RECT 157.920 130.500 158.960 130.800 ;
        RECT 159.120 130.760 159.440 131.090 ;
        RECT 154.590 130.360 158.960 130.500 ;
        RECT 154.590 130.340 157.970 130.360 ;
        RECT 153.540 129.420 155.600 129.690 ;
        RECT 153.540 127.590 153.910 129.420 ;
        RECT 154.160 128.960 154.420 128.990 ;
        RECT 154.160 128.670 154.440 128.960 ;
        RECT 154.600 128.870 155.600 129.420 ;
        RECT 156.470 128.990 157.200 130.340 ;
        RECT 159.690 129.760 160.040 131.590 ;
        RECT 157.920 129.490 160.040 129.760 ;
        RECT 154.600 128.700 155.600 128.710 ;
        RECT 154.160 128.650 154.420 128.670 ;
        RECT 154.590 128.490 155.600 128.700 ;
        RECT 155.740 128.660 157.770 128.990 ;
        RECT 157.930 128.960 158.960 129.490 ;
        RECT 157.945 128.930 158.945 128.960 ;
        RECT 157.945 128.700 158.945 128.720 ;
        RECT 154.590 128.400 155.740 128.490 ;
        RECT 157.920 128.400 158.960 128.700 ;
        RECT 159.120 128.660 159.440 128.990 ;
        RECT 154.590 128.260 158.960 128.400 ;
        RECT 154.590 128.240 157.970 128.260 ;
        RECT 153.540 127.320 155.600 127.590 ;
        RECT 153.540 125.490 153.910 127.320 ;
        RECT 154.160 126.860 154.420 126.890 ;
        RECT 154.160 126.570 154.440 126.860 ;
        RECT 154.600 126.770 155.600 127.320 ;
        RECT 156.470 126.890 157.200 128.240 ;
        RECT 159.690 127.660 160.040 129.490 ;
        RECT 157.920 127.390 160.040 127.660 ;
        RECT 154.600 126.600 155.600 126.610 ;
        RECT 154.160 126.550 154.420 126.570 ;
        RECT 154.590 126.390 155.600 126.600 ;
        RECT 155.740 126.560 157.770 126.890 ;
        RECT 157.930 126.860 158.960 127.390 ;
        RECT 157.945 126.830 158.945 126.860 ;
        RECT 157.945 126.600 158.945 126.620 ;
        RECT 154.590 126.300 155.740 126.390 ;
        RECT 157.920 126.300 158.960 126.600 ;
        RECT 159.120 126.560 159.440 126.890 ;
        RECT 154.590 126.160 158.960 126.300 ;
        RECT 154.590 126.140 157.970 126.160 ;
        RECT 153.540 125.220 155.600 125.490 ;
        RECT 153.540 123.390 153.910 125.220 ;
        RECT 154.160 124.760 154.420 124.790 ;
        RECT 154.160 124.470 154.440 124.760 ;
        RECT 154.600 124.670 155.600 125.220 ;
        RECT 156.470 124.790 157.200 126.140 ;
        RECT 159.690 125.560 160.040 127.390 ;
        RECT 157.920 125.290 160.040 125.560 ;
        RECT 154.600 124.500 155.600 124.510 ;
        RECT 154.160 124.450 154.420 124.470 ;
        RECT 154.590 124.290 155.600 124.500 ;
        RECT 155.740 124.460 157.770 124.790 ;
        RECT 157.930 124.760 158.960 125.290 ;
        RECT 157.945 124.730 158.945 124.760 ;
        RECT 157.945 124.500 158.945 124.520 ;
        RECT 154.590 124.200 155.740 124.290 ;
        RECT 157.920 124.200 158.960 124.500 ;
        RECT 159.120 124.460 159.440 124.790 ;
        RECT 154.590 124.060 158.960 124.200 ;
        RECT 154.590 124.040 157.970 124.060 ;
        RECT 153.540 123.120 155.600 123.390 ;
        RECT 153.540 121.290 153.910 123.120 ;
        RECT 154.160 122.660 154.420 122.690 ;
        RECT 154.160 122.370 154.440 122.660 ;
        RECT 154.600 122.570 155.600 123.120 ;
        RECT 156.470 122.690 157.200 124.040 ;
        RECT 159.690 123.460 160.040 125.290 ;
        RECT 157.920 123.190 160.040 123.460 ;
        RECT 154.600 122.400 155.600 122.410 ;
        RECT 154.160 122.350 154.420 122.370 ;
        RECT 154.590 122.190 155.600 122.400 ;
        RECT 155.740 122.360 157.770 122.690 ;
        RECT 157.930 122.660 158.960 123.190 ;
        RECT 157.945 122.630 158.945 122.660 ;
        RECT 157.945 122.400 158.945 122.420 ;
        RECT 154.590 122.100 155.740 122.190 ;
        RECT 157.920 122.100 158.960 122.400 ;
        RECT 159.120 122.360 159.440 122.690 ;
        RECT 154.590 121.960 158.960 122.100 ;
        RECT 154.590 121.940 157.970 121.960 ;
        RECT 153.540 121.020 155.600 121.290 ;
        RECT 153.540 119.190 153.910 121.020 ;
        RECT 154.160 120.560 154.420 120.590 ;
        RECT 154.160 120.270 154.440 120.560 ;
        RECT 154.600 120.470 155.600 121.020 ;
        RECT 156.470 120.590 157.200 121.940 ;
        RECT 159.690 121.360 160.040 123.190 ;
        RECT 157.920 121.090 160.040 121.360 ;
        RECT 154.600 120.300 155.600 120.310 ;
        RECT 154.160 120.250 154.420 120.270 ;
        RECT 154.590 120.090 155.600 120.300 ;
        RECT 155.740 120.260 157.770 120.590 ;
        RECT 157.930 120.560 158.960 121.090 ;
        RECT 157.945 120.530 158.945 120.560 ;
        RECT 157.945 120.300 158.945 120.320 ;
        RECT 154.590 120.000 155.740 120.090 ;
        RECT 157.920 120.000 158.960 120.300 ;
        RECT 159.120 120.260 159.440 120.590 ;
        RECT 154.590 119.860 158.960 120.000 ;
        RECT 154.590 119.840 157.970 119.860 ;
        RECT 153.540 118.920 155.600 119.190 ;
        RECT 153.540 117.090 153.910 118.920 ;
        RECT 154.160 118.460 154.420 118.490 ;
        RECT 154.160 118.170 154.440 118.460 ;
        RECT 154.600 118.370 155.600 118.920 ;
        RECT 156.470 118.490 157.200 119.840 ;
        RECT 159.690 119.260 160.040 121.090 ;
        RECT 157.920 118.990 160.040 119.260 ;
        RECT 154.600 118.200 155.600 118.210 ;
        RECT 154.160 118.150 154.420 118.170 ;
        RECT 154.590 117.990 155.600 118.200 ;
        RECT 155.740 118.160 157.770 118.490 ;
        RECT 157.930 118.460 158.960 118.990 ;
        RECT 157.945 118.430 158.945 118.460 ;
        RECT 157.945 118.200 158.945 118.220 ;
        RECT 154.590 117.900 155.740 117.990 ;
        RECT 157.920 117.900 158.960 118.200 ;
        RECT 159.120 118.160 159.440 118.490 ;
        RECT 154.590 117.760 158.960 117.900 ;
        RECT 154.590 117.740 157.970 117.760 ;
        RECT 153.540 116.820 155.600 117.090 ;
        RECT 153.540 114.990 153.910 116.820 ;
        RECT 154.160 116.360 154.420 116.390 ;
        RECT 154.160 116.070 154.440 116.360 ;
        RECT 154.600 116.270 155.600 116.820 ;
        RECT 156.470 116.390 157.200 117.740 ;
        RECT 159.690 117.160 160.040 118.990 ;
        RECT 157.920 116.890 160.040 117.160 ;
        RECT 154.600 116.100 155.600 116.110 ;
        RECT 154.160 116.050 154.420 116.070 ;
        RECT 154.590 115.890 155.600 116.100 ;
        RECT 155.740 116.060 157.770 116.390 ;
        RECT 157.930 116.360 158.960 116.890 ;
        RECT 157.945 116.330 158.945 116.360 ;
        RECT 157.945 116.100 158.945 116.120 ;
        RECT 154.590 115.800 155.740 115.890 ;
        RECT 157.920 115.800 158.960 116.100 ;
        RECT 159.120 116.060 159.440 116.390 ;
        RECT 154.590 115.660 158.960 115.800 ;
        RECT 154.590 115.640 157.970 115.660 ;
        RECT 153.540 114.720 155.600 114.990 ;
        RECT 153.540 112.890 153.910 114.720 ;
        RECT 154.160 114.260 154.420 114.290 ;
        RECT 154.160 113.970 154.440 114.260 ;
        RECT 154.600 114.170 155.600 114.720 ;
        RECT 156.470 114.290 157.200 115.640 ;
        RECT 159.690 115.060 160.040 116.890 ;
        RECT 157.920 114.790 160.040 115.060 ;
        RECT 154.600 114.000 155.600 114.010 ;
        RECT 154.160 113.950 154.420 113.970 ;
        RECT 154.590 113.790 155.600 114.000 ;
        RECT 155.740 113.960 157.770 114.290 ;
        RECT 157.930 114.260 158.960 114.790 ;
        RECT 157.945 114.230 158.945 114.260 ;
        RECT 157.945 114.000 158.945 114.020 ;
        RECT 154.590 113.700 155.740 113.790 ;
        RECT 157.920 113.700 158.960 114.000 ;
        RECT 159.120 113.960 159.440 114.290 ;
        RECT 154.590 113.560 158.960 113.700 ;
        RECT 154.590 113.540 157.970 113.560 ;
        RECT 153.540 112.620 155.600 112.890 ;
        RECT 153.540 110.790 153.910 112.620 ;
        RECT 154.160 112.160 154.420 112.190 ;
        RECT 154.160 111.870 154.440 112.160 ;
        RECT 154.600 112.070 155.600 112.620 ;
        RECT 156.470 112.190 157.200 113.540 ;
        RECT 159.690 112.960 160.040 114.790 ;
        RECT 157.920 112.690 160.040 112.960 ;
        RECT 154.600 111.900 155.600 111.910 ;
        RECT 154.160 111.850 154.420 111.870 ;
        RECT 154.590 111.690 155.600 111.900 ;
        RECT 155.740 111.860 157.770 112.190 ;
        RECT 157.930 112.160 158.960 112.690 ;
        RECT 157.945 112.130 158.945 112.160 ;
        RECT 157.945 111.900 158.945 111.920 ;
        RECT 154.590 111.600 155.740 111.690 ;
        RECT 157.920 111.600 158.960 111.900 ;
        RECT 159.120 111.860 159.440 112.190 ;
        RECT 154.590 111.460 158.960 111.600 ;
        RECT 154.590 111.440 157.970 111.460 ;
        RECT 153.540 110.520 155.600 110.790 ;
        RECT 153.540 108.690 153.910 110.520 ;
        RECT 154.160 110.060 154.420 110.090 ;
        RECT 154.160 109.770 154.440 110.060 ;
        RECT 154.600 109.970 155.600 110.520 ;
        RECT 156.470 110.090 157.200 111.440 ;
        RECT 159.690 110.860 160.040 112.690 ;
        RECT 157.920 110.590 160.040 110.860 ;
        RECT 154.600 109.800 155.600 109.810 ;
        RECT 154.160 109.750 154.420 109.770 ;
        RECT 154.590 109.590 155.600 109.800 ;
        RECT 155.740 109.760 157.770 110.090 ;
        RECT 157.930 110.060 158.960 110.590 ;
        RECT 157.945 110.030 158.945 110.060 ;
        RECT 157.945 109.800 158.945 109.820 ;
        RECT 154.590 109.500 155.740 109.590 ;
        RECT 157.920 109.500 158.960 109.800 ;
        RECT 159.120 109.760 159.440 110.090 ;
        RECT 154.590 109.360 158.960 109.500 ;
        RECT 154.590 109.340 157.970 109.360 ;
        RECT 153.540 108.420 155.600 108.690 ;
        RECT 153.540 106.590 153.910 108.420 ;
        RECT 154.160 107.960 154.420 107.990 ;
        RECT 154.160 107.670 154.440 107.960 ;
        RECT 154.600 107.870 155.600 108.420 ;
        RECT 156.470 107.990 157.200 109.340 ;
        RECT 159.690 108.760 160.040 110.590 ;
        RECT 157.920 108.490 160.040 108.760 ;
        RECT 154.600 107.700 155.600 107.710 ;
        RECT 154.160 107.650 154.420 107.670 ;
        RECT 154.590 107.490 155.600 107.700 ;
        RECT 155.740 107.660 157.770 107.990 ;
        RECT 157.930 107.960 158.960 108.490 ;
        RECT 157.945 107.930 158.945 107.960 ;
        RECT 157.945 107.700 158.945 107.720 ;
        RECT 154.590 107.400 155.740 107.490 ;
        RECT 157.920 107.400 158.960 107.700 ;
        RECT 159.120 107.660 159.440 107.990 ;
        RECT 154.590 107.260 158.960 107.400 ;
        RECT 154.590 107.240 157.970 107.260 ;
        RECT 153.540 106.320 155.600 106.590 ;
        RECT 153.540 104.490 153.910 106.320 ;
        RECT 154.160 105.860 154.420 105.890 ;
        RECT 154.160 105.570 154.440 105.860 ;
        RECT 154.600 105.770 155.600 106.320 ;
        RECT 156.470 105.890 157.200 107.240 ;
        RECT 159.690 106.660 160.040 108.490 ;
        RECT 157.920 106.390 160.040 106.660 ;
        RECT 154.600 105.600 155.600 105.610 ;
        RECT 154.160 105.550 154.420 105.570 ;
        RECT 154.590 105.390 155.600 105.600 ;
        RECT 155.740 105.560 157.770 105.890 ;
        RECT 157.930 105.860 158.960 106.390 ;
        RECT 157.945 105.830 158.945 105.860 ;
        RECT 157.945 105.600 158.945 105.620 ;
        RECT 154.590 105.300 155.740 105.390 ;
        RECT 157.920 105.300 158.960 105.600 ;
        RECT 159.120 105.560 159.440 105.890 ;
        RECT 154.590 105.160 158.960 105.300 ;
        RECT 154.590 105.140 157.970 105.160 ;
        RECT 153.540 104.220 155.600 104.490 ;
        RECT 153.540 102.390 153.910 104.220 ;
        RECT 154.160 103.760 154.420 103.790 ;
        RECT 154.160 103.470 154.440 103.760 ;
        RECT 154.600 103.670 155.600 104.220 ;
        RECT 156.470 103.790 157.200 105.140 ;
        RECT 159.690 104.560 160.040 106.390 ;
        RECT 157.920 104.290 160.040 104.560 ;
        RECT 154.600 103.500 155.600 103.510 ;
        RECT 154.160 103.450 154.420 103.470 ;
        RECT 154.590 103.290 155.600 103.500 ;
        RECT 155.740 103.460 157.770 103.790 ;
        RECT 157.930 103.760 158.960 104.290 ;
        RECT 157.945 103.730 158.945 103.760 ;
        RECT 157.945 103.500 158.945 103.520 ;
        RECT 154.590 103.200 155.740 103.290 ;
        RECT 157.920 103.200 158.960 103.500 ;
        RECT 159.120 103.460 159.440 103.790 ;
        RECT 154.590 103.060 158.960 103.200 ;
        RECT 154.590 103.040 157.970 103.060 ;
        RECT 153.540 102.120 155.600 102.390 ;
        RECT 153.540 100.290 153.910 102.120 ;
        RECT 154.160 101.660 154.420 101.690 ;
        RECT 154.160 101.370 154.440 101.660 ;
        RECT 154.600 101.570 155.600 102.120 ;
        RECT 156.470 101.690 157.200 103.040 ;
        RECT 159.690 102.460 160.040 104.290 ;
        RECT 157.920 102.190 160.040 102.460 ;
        RECT 154.600 101.400 155.600 101.410 ;
        RECT 154.160 101.350 154.420 101.370 ;
        RECT 154.590 101.190 155.600 101.400 ;
        RECT 155.740 101.360 157.770 101.690 ;
        RECT 157.930 101.660 158.960 102.190 ;
        RECT 157.945 101.630 158.945 101.660 ;
        RECT 157.945 101.400 158.945 101.420 ;
        RECT 154.590 101.100 155.740 101.190 ;
        RECT 157.920 101.100 158.960 101.400 ;
        RECT 159.120 101.360 159.440 101.690 ;
        RECT 154.590 100.960 158.960 101.100 ;
        RECT 154.590 100.940 157.970 100.960 ;
        RECT 153.540 100.020 155.600 100.290 ;
        RECT 153.540 98.190 153.910 100.020 ;
        RECT 154.160 99.560 154.420 99.590 ;
        RECT 154.160 99.270 154.440 99.560 ;
        RECT 154.600 99.470 155.600 100.020 ;
        RECT 156.470 99.590 157.200 100.940 ;
        RECT 159.690 100.360 160.040 102.190 ;
        RECT 157.920 100.090 160.040 100.360 ;
        RECT 154.600 99.300 155.600 99.310 ;
        RECT 154.160 99.250 154.420 99.270 ;
        RECT 154.590 99.090 155.600 99.300 ;
        RECT 155.740 99.260 157.770 99.590 ;
        RECT 157.930 99.560 158.960 100.090 ;
        RECT 157.945 99.530 158.945 99.560 ;
        RECT 157.945 99.300 158.945 99.320 ;
        RECT 154.590 99.000 155.740 99.090 ;
        RECT 157.920 99.000 158.960 99.300 ;
        RECT 159.120 99.260 159.440 99.590 ;
        RECT 154.590 98.860 158.960 99.000 ;
        RECT 154.590 98.840 157.970 98.860 ;
        RECT 153.540 97.920 155.600 98.190 ;
        RECT 153.540 96.090 153.910 97.920 ;
        RECT 154.160 97.460 154.420 97.490 ;
        RECT 154.160 97.170 154.440 97.460 ;
        RECT 154.600 97.370 155.600 97.920 ;
        RECT 156.470 97.490 157.200 98.840 ;
        RECT 159.690 98.260 160.040 100.090 ;
        RECT 157.920 97.990 160.040 98.260 ;
        RECT 154.600 97.200 155.600 97.210 ;
        RECT 154.160 97.150 154.420 97.170 ;
        RECT 154.590 96.990 155.600 97.200 ;
        RECT 155.740 97.160 157.770 97.490 ;
        RECT 157.930 97.460 158.960 97.990 ;
        RECT 157.945 97.430 158.945 97.460 ;
        RECT 157.945 97.200 158.945 97.220 ;
        RECT 154.590 96.900 155.740 96.990 ;
        RECT 157.920 96.900 158.960 97.200 ;
        RECT 159.120 97.160 159.440 97.490 ;
        RECT 154.590 96.760 158.960 96.900 ;
        RECT 154.590 96.740 157.970 96.760 ;
        RECT 153.540 95.820 155.600 96.090 ;
        RECT 153.540 93.990 153.910 95.820 ;
        RECT 154.160 95.360 154.420 95.390 ;
        RECT 154.160 95.070 154.440 95.360 ;
        RECT 154.600 95.270 155.600 95.820 ;
        RECT 156.470 95.390 157.200 96.740 ;
        RECT 159.690 96.160 160.040 97.990 ;
        RECT 157.920 95.890 160.040 96.160 ;
        RECT 154.600 95.100 155.600 95.110 ;
        RECT 154.160 95.050 154.420 95.070 ;
        RECT 154.590 94.890 155.600 95.100 ;
        RECT 155.740 95.060 157.770 95.390 ;
        RECT 157.930 95.360 158.960 95.890 ;
        RECT 157.945 95.330 158.945 95.360 ;
        RECT 157.945 95.100 158.945 95.120 ;
        RECT 154.590 94.800 155.740 94.890 ;
        RECT 157.920 94.800 158.960 95.100 ;
        RECT 159.120 95.060 159.440 95.390 ;
        RECT 154.590 94.660 158.960 94.800 ;
        RECT 154.590 94.640 157.970 94.660 ;
        RECT 153.540 93.720 155.600 93.990 ;
        RECT 153.540 91.890 153.910 93.720 ;
        RECT 154.160 93.260 154.420 93.290 ;
        RECT 154.160 92.970 154.440 93.260 ;
        RECT 154.600 93.170 155.600 93.720 ;
        RECT 156.470 93.290 157.200 94.640 ;
        RECT 159.690 94.060 160.040 95.890 ;
        RECT 157.920 93.790 160.040 94.060 ;
        RECT 154.600 93.000 155.600 93.010 ;
        RECT 154.160 92.950 154.420 92.970 ;
        RECT 154.590 92.790 155.600 93.000 ;
        RECT 155.740 92.960 157.770 93.290 ;
        RECT 157.930 93.260 158.960 93.790 ;
        RECT 157.945 93.230 158.945 93.260 ;
        RECT 157.945 93.000 158.945 93.020 ;
        RECT 154.590 92.700 155.740 92.790 ;
        RECT 157.920 92.700 158.960 93.000 ;
        RECT 159.120 92.960 159.440 93.290 ;
        RECT 154.590 92.560 158.960 92.700 ;
        RECT 154.590 92.540 157.970 92.560 ;
        RECT 153.540 91.620 155.600 91.890 ;
        RECT 153.540 89.790 153.910 91.620 ;
        RECT 154.160 91.160 154.420 91.190 ;
        RECT 154.160 90.870 154.440 91.160 ;
        RECT 154.600 91.070 155.600 91.620 ;
        RECT 156.470 91.190 157.200 92.540 ;
        RECT 159.690 91.960 160.040 93.790 ;
        RECT 157.920 91.690 160.040 91.960 ;
        RECT 154.600 90.900 155.600 90.910 ;
        RECT 154.160 90.850 154.420 90.870 ;
        RECT 154.590 90.690 155.600 90.900 ;
        RECT 155.740 90.860 157.770 91.190 ;
        RECT 157.930 91.160 158.960 91.690 ;
        RECT 157.945 91.130 158.945 91.160 ;
        RECT 157.945 90.900 158.945 90.920 ;
        RECT 154.590 90.600 155.740 90.690 ;
        RECT 157.920 90.600 158.960 90.900 ;
        RECT 159.120 90.860 159.440 91.190 ;
        RECT 154.590 90.460 158.960 90.600 ;
        RECT 154.590 90.440 157.970 90.460 ;
        RECT 153.540 89.520 155.600 89.790 ;
        RECT 153.540 87.690 153.910 89.520 ;
        RECT 154.160 89.060 154.420 89.090 ;
        RECT 154.160 88.770 154.440 89.060 ;
        RECT 154.600 88.970 155.600 89.520 ;
        RECT 156.470 89.090 157.200 90.440 ;
        RECT 159.690 89.860 160.040 91.690 ;
        RECT 157.920 89.590 160.040 89.860 ;
        RECT 154.600 88.800 155.600 88.810 ;
        RECT 154.160 88.750 154.420 88.770 ;
        RECT 154.590 88.590 155.600 88.800 ;
        RECT 155.740 88.760 157.770 89.090 ;
        RECT 157.930 89.060 158.960 89.590 ;
        RECT 157.945 89.030 158.945 89.060 ;
        RECT 157.945 88.800 158.945 88.820 ;
        RECT 154.590 88.500 155.740 88.590 ;
        RECT 157.920 88.500 158.960 88.800 ;
        RECT 159.120 88.760 159.440 89.090 ;
        RECT 154.590 88.360 158.960 88.500 ;
        RECT 154.590 88.340 157.970 88.360 ;
        RECT 153.540 87.420 155.600 87.690 ;
        RECT 153.540 85.590 153.910 87.420 ;
        RECT 154.160 86.960 154.420 86.990 ;
        RECT 154.160 86.670 154.440 86.960 ;
        RECT 154.600 86.870 155.600 87.420 ;
        RECT 156.470 86.990 157.200 88.340 ;
        RECT 159.690 87.760 160.040 89.590 ;
        RECT 157.920 87.490 160.040 87.760 ;
        RECT 154.600 86.700 155.600 86.710 ;
        RECT 154.160 86.650 154.420 86.670 ;
        RECT 154.590 86.490 155.600 86.700 ;
        RECT 155.740 86.660 157.770 86.990 ;
        RECT 157.930 86.960 158.960 87.490 ;
        RECT 157.945 86.930 158.945 86.960 ;
        RECT 157.945 86.700 158.945 86.720 ;
        RECT 154.590 86.400 155.740 86.490 ;
        RECT 157.920 86.400 158.960 86.700 ;
        RECT 159.120 86.660 159.440 86.990 ;
        RECT 154.590 86.260 158.960 86.400 ;
        RECT 154.590 86.240 157.970 86.260 ;
        RECT 153.540 85.320 155.600 85.590 ;
        RECT 153.540 83.490 153.910 85.320 ;
        RECT 154.160 84.860 154.420 84.890 ;
        RECT 154.160 84.570 154.440 84.860 ;
        RECT 154.600 84.770 155.600 85.320 ;
        RECT 156.470 84.890 157.200 86.240 ;
        RECT 159.690 85.660 160.040 87.490 ;
        RECT 157.920 85.390 160.040 85.660 ;
        RECT 154.600 84.600 155.600 84.610 ;
        RECT 154.160 84.550 154.420 84.570 ;
        RECT 154.590 84.390 155.600 84.600 ;
        RECT 155.740 84.560 157.770 84.890 ;
        RECT 157.930 84.860 158.960 85.390 ;
        RECT 157.945 84.830 158.945 84.860 ;
        RECT 157.945 84.600 158.945 84.620 ;
        RECT 154.590 84.300 155.740 84.390 ;
        RECT 157.920 84.300 158.960 84.600 ;
        RECT 159.120 84.560 159.440 84.890 ;
        RECT 154.590 84.160 158.960 84.300 ;
        RECT 154.590 84.140 157.970 84.160 ;
        RECT 153.540 83.220 155.600 83.490 ;
        RECT 153.540 81.390 153.910 83.220 ;
        RECT 154.160 82.760 154.420 82.790 ;
        RECT 154.160 82.470 154.440 82.760 ;
        RECT 154.600 82.670 155.600 83.220 ;
        RECT 156.470 82.790 157.200 84.140 ;
        RECT 159.690 83.560 160.040 85.390 ;
        RECT 157.920 83.290 160.040 83.560 ;
        RECT 154.600 82.500 155.600 82.510 ;
        RECT 154.160 82.450 154.420 82.470 ;
        RECT 154.590 82.290 155.600 82.500 ;
        RECT 155.740 82.460 157.770 82.790 ;
        RECT 157.930 82.760 158.960 83.290 ;
        RECT 157.945 82.730 158.945 82.760 ;
        RECT 157.945 82.500 158.945 82.520 ;
        RECT 154.590 82.200 155.740 82.290 ;
        RECT 157.920 82.200 158.960 82.500 ;
        RECT 159.120 82.460 159.440 82.790 ;
        RECT 154.590 82.060 158.960 82.200 ;
        RECT 154.590 82.040 157.970 82.060 ;
        RECT 153.540 81.120 155.600 81.390 ;
        RECT 153.540 79.290 153.910 81.120 ;
        RECT 154.160 80.660 154.420 80.690 ;
        RECT 154.160 80.370 154.440 80.660 ;
        RECT 154.600 80.570 155.600 81.120 ;
        RECT 156.470 80.690 157.200 82.040 ;
        RECT 159.690 81.460 160.040 83.290 ;
        RECT 157.920 81.190 160.040 81.460 ;
        RECT 154.600 80.400 155.600 80.410 ;
        RECT 154.160 80.350 154.420 80.370 ;
        RECT 154.590 80.190 155.600 80.400 ;
        RECT 155.740 80.360 157.770 80.690 ;
        RECT 157.930 80.660 158.960 81.190 ;
        RECT 157.945 80.630 158.945 80.660 ;
        RECT 157.945 80.400 158.945 80.420 ;
        RECT 154.590 80.100 155.740 80.190 ;
        RECT 157.920 80.100 158.960 80.400 ;
        RECT 159.120 80.360 159.440 80.690 ;
        RECT 154.590 79.960 158.960 80.100 ;
        RECT 154.590 79.940 157.970 79.960 ;
        RECT 153.540 79.020 155.600 79.290 ;
        RECT 153.540 77.190 153.910 79.020 ;
        RECT 154.160 78.560 154.420 78.590 ;
        RECT 154.160 78.270 154.440 78.560 ;
        RECT 154.600 78.470 155.600 79.020 ;
        RECT 156.470 78.590 157.200 79.940 ;
        RECT 159.690 79.360 160.040 81.190 ;
        RECT 157.920 79.090 160.040 79.360 ;
        RECT 154.600 78.300 155.600 78.310 ;
        RECT 154.160 78.250 154.420 78.270 ;
        RECT 154.590 78.090 155.600 78.300 ;
        RECT 155.740 78.260 157.770 78.590 ;
        RECT 157.930 78.560 158.960 79.090 ;
        RECT 157.945 78.530 158.945 78.560 ;
        RECT 157.945 78.300 158.945 78.320 ;
        RECT 154.590 78.000 155.740 78.090 ;
        RECT 157.920 78.000 158.960 78.300 ;
        RECT 159.120 78.260 159.440 78.590 ;
        RECT 154.590 77.860 158.960 78.000 ;
        RECT 154.590 77.840 157.970 77.860 ;
        RECT 153.540 76.920 155.600 77.190 ;
        RECT 153.540 75.090 153.910 76.920 ;
        RECT 154.160 76.460 154.420 76.490 ;
        RECT 154.160 76.170 154.440 76.460 ;
        RECT 154.600 76.370 155.600 76.920 ;
        RECT 156.470 76.490 157.200 77.840 ;
        RECT 159.690 77.260 160.040 79.090 ;
        RECT 157.920 76.990 160.040 77.260 ;
        RECT 154.600 76.200 155.600 76.210 ;
        RECT 154.160 76.150 154.420 76.170 ;
        RECT 154.590 75.990 155.600 76.200 ;
        RECT 155.740 76.160 157.770 76.490 ;
        RECT 157.930 76.460 158.960 76.990 ;
        RECT 157.945 76.430 158.945 76.460 ;
        RECT 157.945 76.200 158.945 76.220 ;
        RECT 154.590 75.900 155.740 75.990 ;
        RECT 157.920 75.900 158.960 76.200 ;
        RECT 159.120 76.160 159.440 76.490 ;
        RECT 154.590 75.760 158.960 75.900 ;
        RECT 154.590 75.740 157.970 75.760 ;
        RECT 153.540 74.820 155.600 75.090 ;
        RECT 153.540 72.990 153.910 74.820 ;
        RECT 154.160 74.360 154.420 74.390 ;
        RECT 154.160 74.070 154.440 74.360 ;
        RECT 154.600 74.270 155.600 74.820 ;
        RECT 156.470 74.390 157.200 75.740 ;
        RECT 159.690 75.160 160.040 76.990 ;
        RECT 157.920 74.890 160.040 75.160 ;
        RECT 154.600 74.100 155.600 74.110 ;
        RECT 154.160 74.050 154.420 74.070 ;
        RECT 154.590 73.890 155.600 74.100 ;
        RECT 155.740 74.060 157.770 74.390 ;
        RECT 157.930 74.360 158.960 74.890 ;
        RECT 157.945 74.330 158.945 74.360 ;
        RECT 157.945 74.100 158.945 74.120 ;
        RECT 154.590 73.800 155.740 73.890 ;
        RECT 157.920 73.800 158.960 74.100 ;
        RECT 159.120 74.060 159.440 74.390 ;
        RECT 154.590 73.660 158.960 73.800 ;
        RECT 154.590 73.640 157.970 73.660 ;
        RECT 153.540 72.720 155.600 72.990 ;
        RECT 153.540 70.890 153.910 72.720 ;
        RECT 154.160 72.260 154.420 72.290 ;
        RECT 154.160 71.970 154.440 72.260 ;
        RECT 154.600 72.170 155.600 72.720 ;
        RECT 156.470 72.290 157.200 73.640 ;
        RECT 159.690 73.060 160.040 74.890 ;
        RECT 157.920 72.790 160.040 73.060 ;
        RECT 154.600 72.000 155.600 72.010 ;
        RECT 154.160 71.950 154.420 71.970 ;
        RECT 154.590 71.790 155.600 72.000 ;
        RECT 155.740 71.960 157.770 72.290 ;
        RECT 157.930 72.260 158.960 72.790 ;
        RECT 157.945 72.230 158.945 72.260 ;
        RECT 157.945 72.000 158.945 72.020 ;
        RECT 154.590 71.700 155.740 71.790 ;
        RECT 157.920 71.700 158.960 72.000 ;
        RECT 159.120 71.960 159.440 72.290 ;
        RECT 154.590 71.560 158.960 71.700 ;
        RECT 154.590 71.540 157.970 71.560 ;
        RECT 153.540 70.620 155.600 70.890 ;
        RECT 153.540 68.790 153.910 70.620 ;
        RECT 154.160 70.160 154.420 70.190 ;
        RECT 154.160 69.870 154.440 70.160 ;
        RECT 154.600 70.070 155.600 70.620 ;
        RECT 156.470 70.190 157.200 71.540 ;
        RECT 159.690 70.960 160.040 72.790 ;
        RECT 157.920 70.690 160.040 70.960 ;
        RECT 154.600 69.900 155.600 69.910 ;
        RECT 154.160 69.850 154.420 69.870 ;
        RECT 154.590 69.690 155.600 69.900 ;
        RECT 155.740 69.860 157.770 70.190 ;
        RECT 157.930 70.160 158.960 70.690 ;
        RECT 157.945 70.130 158.945 70.160 ;
        RECT 157.945 69.900 158.945 69.920 ;
        RECT 154.590 69.600 155.740 69.690 ;
        RECT 157.920 69.600 158.960 69.900 ;
        RECT 159.120 69.860 159.440 70.190 ;
        RECT 154.590 69.460 158.960 69.600 ;
        RECT 154.590 69.440 157.970 69.460 ;
        RECT 153.540 68.520 155.600 68.790 ;
        RECT 153.540 66.690 153.910 68.520 ;
        RECT 154.160 68.060 154.420 68.090 ;
        RECT 154.160 67.770 154.440 68.060 ;
        RECT 154.600 67.970 155.600 68.520 ;
        RECT 156.470 68.090 157.200 69.440 ;
        RECT 159.690 68.860 160.040 70.690 ;
        RECT 157.920 68.590 160.040 68.860 ;
        RECT 154.600 67.800 155.600 67.810 ;
        RECT 154.160 67.750 154.420 67.770 ;
        RECT 154.590 67.590 155.600 67.800 ;
        RECT 155.740 67.760 157.770 68.090 ;
        RECT 157.930 68.060 158.960 68.590 ;
        RECT 157.945 68.030 158.945 68.060 ;
        RECT 157.945 67.800 158.945 67.820 ;
        RECT 154.590 67.500 155.740 67.590 ;
        RECT 157.920 67.500 158.960 67.800 ;
        RECT 159.120 67.760 159.440 68.090 ;
        RECT 154.590 67.360 158.960 67.500 ;
        RECT 154.590 67.340 157.970 67.360 ;
        RECT 153.540 66.420 155.600 66.690 ;
        RECT 153.540 64.590 153.910 66.420 ;
        RECT 154.160 65.960 154.420 65.990 ;
        RECT 154.160 65.670 154.440 65.960 ;
        RECT 154.600 65.870 155.600 66.420 ;
        RECT 156.470 65.990 157.200 67.340 ;
        RECT 159.690 66.760 160.040 68.590 ;
        RECT 157.920 66.490 160.040 66.760 ;
        RECT 154.600 65.700 155.600 65.710 ;
        RECT 154.160 65.650 154.420 65.670 ;
        RECT 154.590 65.490 155.600 65.700 ;
        RECT 155.740 65.660 157.770 65.990 ;
        RECT 157.930 65.960 158.960 66.490 ;
        RECT 157.945 65.930 158.945 65.960 ;
        RECT 157.945 65.700 158.945 65.720 ;
        RECT 154.590 65.400 155.740 65.490 ;
        RECT 157.920 65.400 158.960 65.700 ;
        RECT 159.120 65.660 159.440 65.990 ;
        RECT 154.590 65.260 158.960 65.400 ;
        RECT 154.590 65.240 157.970 65.260 ;
        RECT 153.540 64.320 155.600 64.590 ;
        RECT 153.540 62.490 153.910 64.320 ;
        RECT 154.160 63.860 154.420 63.890 ;
        RECT 154.160 63.570 154.440 63.860 ;
        RECT 154.600 63.770 155.600 64.320 ;
        RECT 156.470 63.890 157.200 65.240 ;
        RECT 159.690 64.660 160.040 66.490 ;
        RECT 157.920 64.390 160.040 64.660 ;
        RECT 154.600 63.600 155.600 63.610 ;
        RECT 154.160 63.550 154.420 63.570 ;
        RECT 154.590 63.390 155.600 63.600 ;
        RECT 155.740 63.560 157.770 63.890 ;
        RECT 157.930 63.860 158.960 64.390 ;
        RECT 157.945 63.830 158.945 63.860 ;
        RECT 157.945 63.600 158.945 63.620 ;
        RECT 154.590 63.300 155.740 63.390 ;
        RECT 157.920 63.300 158.960 63.600 ;
        RECT 159.120 63.560 159.440 63.890 ;
        RECT 154.590 63.160 158.960 63.300 ;
        RECT 154.590 63.140 157.970 63.160 ;
        RECT 153.540 62.220 155.600 62.490 ;
        RECT 153.540 60.390 153.910 62.220 ;
        RECT 154.160 61.760 154.420 61.790 ;
        RECT 154.160 61.470 154.440 61.760 ;
        RECT 154.600 61.670 155.600 62.220 ;
        RECT 156.470 61.790 157.200 63.140 ;
        RECT 159.690 62.560 160.040 64.390 ;
        RECT 157.920 62.290 160.040 62.560 ;
        RECT 154.600 61.500 155.600 61.510 ;
        RECT 154.160 61.450 154.420 61.470 ;
        RECT 154.590 61.290 155.600 61.500 ;
        RECT 155.740 61.460 157.770 61.790 ;
        RECT 157.930 61.760 158.960 62.290 ;
        RECT 157.945 61.730 158.945 61.760 ;
        RECT 157.945 61.500 158.945 61.520 ;
        RECT 154.590 61.200 155.740 61.290 ;
        RECT 157.920 61.200 158.960 61.500 ;
        RECT 159.120 61.460 159.440 61.790 ;
        RECT 154.590 61.060 158.960 61.200 ;
        RECT 154.590 61.040 157.970 61.060 ;
        RECT 153.540 60.120 155.600 60.390 ;
        RECT 153.540 58.290 153.910 60.120 ;
        RECT 154.160 59.660 154.420 59.690 ;
        RECT 154.160 59.370 154.440 59.660 ;
        RECT 154.600 59.570 155.600 60.120 ;
        RECT 156.470 59.690 157.200 61.040 ;
        RECT 159.690 60.460 160.040 62.290 ;
        RECT 157.920 60.190 160.040 60.460 ;
        RECT 154.600 59.400 155.600 59.410 ;
        RECT 154.160 59.350 154.420 59.370 ;
        RECT 154.590 59.190 155.600 59.400 ;
        RECT 155.740 59.360 157.770 59.690 ;
        RECT 157.930 59.660 158.960 60.190 ;
        RECT 157.945 59.630 158.945 59.660 ;
        RECT 157.945 59.400 158.945 59.420 ;
        RECT 154.590 59.100 155.740 59.190 ;
        RECT 157.920 59.100 158.960 59.400 ;
        RECT 159.120 59.360 159.440 59.690 ;
        RECT 154.590 58.960 158.960 59.100 ;
        RECT 154.590 58.940 157.970 58.960 ;
        RECT 153.540 58.020 155.600 58.290 ;
        RECT 153.540 56.190 153.910 58.020 ;
        RECT 154.160 57.560 154.420 57.590 ;
        RECT 154.160 57.270 154.440 57.560 ;
        RECT 154.600 57.470 155.600 58.020 ;
        RECT 156.470 57.590 157.200 58.940 ;
        RECT 159.690 58.360 160.040 60.190 ;
        RECT 157.920 58.090 160.040 58.360 ;
        RECT 154.600 57.300 155.600 57.310 ;
        RECT 154.160 57.250 154.420 57.270 ;
        RECT 154.590 57.090 155.600 57.300 ;
        RECT 155.740 57.260 157.770 57.590 ;
        RECT 157.930 57.560 158.960 58.090 ;
        RECT 157.945 57.530 158.945 57.560 ;
        RECT 157.945 57.300 158.945 57.320 ;
        RECT 154.590 57.000 155.740 57.090 ;
        RECT 157.920 57.000 158.960 57.300 ;
        RECT 159.120 57.260 159.440 57.590 ;
        RECT 154.590 56.860 158.960 57.000 ;
        RECT 154.590 56.840 157.970 56.860 ;
        RECT 153.540 55.920 155.600 56.190 ;
        RECT 153.540 54.090 153.910 55.920 ;
        RECT 154.160 55.460 154.420 55.490 ;
        RECT 154.160 55.170 154.440 55.460 ;
        RECT 154.600 55.370 155.600 55.920 ;
        RECT 156.470 55.490 157.200 56.840 ;
        RECT 159.690 56.260 160.040 58.090 ;
        RECT 157.920 55.990 160.040 56.260 ;
        RECT 154.600 55.200 155.600 55.210 ;
        RECT 154.160 55.150 154.420 55.170 ;
        RECT 154.590 54.990 155.600 55.200 ;
        RECT 155.740 55.160 157.770 55.490 ;
        RECT 157.930 55.460 158.960 55.990 ;
        RECT 157.945 55.430 158.945 55.460 ;
        RECT 157.945 55.200 158.945 55.220 ;
        RECT 154.590 54.900 155.740 54.990 ;
        RECT 157.920 54.900 158.960 55.200 ;
        RECT 159.120 55.160 159.440 55.490 ;
        RECT 154.590 54.760 158.960 54.900 ;
        RECT 154.590 54.740 157.970 54.760 ;
        RECT 153.540 53.820 155.600 54.090 ;
        RECT 153.540 51.990 153.910 53.820 ;
        RECT 154.160 53.360 154.420 53.390 ;
        RECT 154.160 53.070 154.440 53.360 ;
        RECT 154.600 53.270 155.600 53.820 ;
        RECT 156.470 53.390 157.200 54.740 ;
        RECT 159.690 54.160 160.040 55.990 ;
        RECT 157.920 53.890 160.040 54.160 ;
        RECT 154.600 53.100 155.600 53.110 ;
        RECT 154.160 53.050 154.420 53.070 ;
        RECT 154.590 52.890 155.600 53.100 ;
        RECT 155.740 53.060 157.770 53.390 ;
        RECT 157.930 53.360 158.960 53.890 ;
        RECT 157.945 53.330 158.945 53.360 ;
        RECT 157.945 53.100 158.945 53.120 ;
        RECT 154.590 52.800 155.740 52.890 ;
        RECT 157.920 52.800 158.960 53.100 ;
        RECT 159.120 53.060 159.440 53.390 ;
        RECT 154.590 52.660 158.960 52.800 ;
        RECT 154.590 52.640 157.970 52.660 ;
        RECT 153.540 51.720 155.600 51.990 ;
        RECT 153.540 49.890 153.910 51.720 ;
        RECT 154.160 51.260 154.420 51.290 ;
        RECT 154.160 50.970 154.440 51.260 ;
        RECT 154.600 51.170 155.600 51.720 ;
        RECT 156.470 51.290 157.200 52.640 ;
        RECT 159.690 52.060 160.040 53.890 ;
        RECT 157.920 51.790 160.040 52.060 ;
        RECT 154.600 51.000 155.600 51.010 ;
        RECT 154.160 50.950 154.420 50.970 ;
        RECT 154.590 50.790 155.600 51.000 ;
        RECT 155.740 50.960 157.770 51.290 ;
        RECT 157.930 51.260 158.960 51.790 ;
        RECT 157.945 51.230 158.945 51.260 ;
        RECT 157.945 51.000 158.945 51.020 ;
        RECT 154.590 50.700 155.740 50.790 ;
        RECT 157.920 50.700 158.960 51.000 ;
        RECT 159.120 50.960 159.440 51.290 ;
        RECT 154.590 50.560 158.960 50.700 ;
        RECT 154.590 50.540 157.970 50.560 ;
        RECT 153.540 49.620 155.600 49.890 ;
        RECT 153.540 47.790 153.910 49.620 ;
        RECT 154.160 49.160 154.420 49.190 ;
        RECT 154.160 48.870 154.440 49.160 ;
        RECT 154.600 49.070 155.600 49.620 ;
        RECT 156.470 49.190 157.200 50.540 ;
        RECT 159.690 49.960 160.040 51.790 ;
        RECT 157.920 49.690 160.040 49.960 ;
        RECT 154.600 48.900 155.600 48.910 ;
        RECT 154.160 48.850 154.420 48.870 ;
        RECT 154.590 48.690 155.600 48.900 ;
        RECT 155.740 48.860 157.770 49.190 ;
        RECT 157.930 49.160 158.960 49.690 ;
        RECT 157.945 49.130 158.945 49.160 ;
        RECT 157.945 48.900 158.945 48.920 ;
        RECT 154.590 48.600 155.740 48.690 ;
        RECT 157.920 48.600 158.960 48.900 ;
        RECT 159.120 48.860 159.440 49.190 ;
        RECT 154.590 48.460 158.960 48.600 ;
        RECT 154.590 48.440 157.970 48.460 ;
        RECT 153.540 47.520 155.600 47.790 ;
        RECT 153.540 45.690 153.910 47.520 ;
        RECT 154.160 47.060 154.420 47.090 ;
        RECT 154.160 46.770 154.440 47.060 ;
        RECT 154.600 46.970 155.600 47.520 ;
        RECT 156.470 47.090 157.200 48.440 ;
        RECT 159.690 47.860 160.040 49.690 ;
        RECT 157.920 47.590 160.040 47.860 ;
        RECT 154.600 46.800 155.600 46.810 ;
        RECT 154.160 46.750 154.420 46.770 ;
        RECT 154.590 46.590 155.600 46.800 ;
        RECT 155.740 46.760 157.770 47.090 ;
        RECT 157.930 47.060 158.960 47.590 ;
        RECT 157.945 47.030 158.945 47.060 ;
        RECT 157.945 46.800 158.945 46.820 ;
        RECT 154.590 46.500 155.740 46.590 ;
        RECT 157.920 46.500 158.960 46.800 ;
        RECT 159.120 46.760 159.440 47.090 ;
        RECT 154.590 46.360 158.960 46.500 ;
        RECT 154.590 46.340 157.970 46.360 ;
        RECT 153.540 45.420 155.600 45.690 ;
        RECT 153.540 43.590 153.910 45.420 ;
        RECT 154.160 44.960 154.420 44.990 ;
        RECT 154.160 44.670 154.440 44.960 ;
        RECT 154.600 44.870 155.600 45.420 ;
        RECT 156.470 44.990 157.200 46.340 ;
        RECT 159.690 45.760 160.040 47.590 ;
        RECT 157.920 45.490 160.040 45.760 ;
        RECT 154.600 44.700 155.600 44.710 ;
        RECT 154.160 44.650 154.420 44.670 ;
        RECT 154.590 44.490 155.600 44.700 ;
        RECT 155.740 44.660 157.770 44.990 ;
        RECT 157.930 44.960 158.960 45.490 ;
        RECT 157.945 44.930 158.945 44.960 ;
        RECT 157.945 44.700 158.945 44.720 ;
        RECT 154.590 44.400 155.740 44.490 ;
        RECT 157.920 44.400 158.960 44.700 ;
        RECT 159.120 44.660 159.440 44.990 ;
        RECT 154.590 44.260 158.960 44.400 ;
        RECT 154.590 44.240 157.970 44.260 ;
        RECT 153.540 43.320 155.600 43.590 ;
        RECT 153.540 41.490 153.910 43.320 ;
        RECT 154.160 42.860 154.420 42.890 ;
        RECT 154.160 42.570 154.440 42.860 ;
        RECT 154.600 42.770 155.600 43.320 ;
        RECT 156.470 42.890 157.200 44.240 ;
        RECT 159.690 43.660 160.040 45.490 ;
        RECT 157.920 43.390 160.040 43.660 ;
        RECT 154.600 42.600 155.600 42.610 ;
        RECT 154.160 42.550 154.420 42.570 ;
        RECT 154.590 42.390 155.600 42.600 ;
        RECT 155.740 42.560 157.770 42.890 ;
        RECT 157.930 42.860 158.960 43.390 ;
        RECT 157.945 42.830 158.945 42.860 ;
        RECT 157.945 42.600 158.945 42.620 ;
        RECT 154.590 42.300 155.740 42.390 ;
        RECT 157.920 42.300 158.960 42.600 ;
        RECT 159.120 42.560 159.440 42.890 ;
        RECT 154.590 42.160 158.960 42.300 ;
        RECT 154.590 42.140 157.970 42.160 ;
        RECT 153.540 41.220 155.600 41.490 ;
        RECT 153.540 39.390 153.910 41.220 ;
        RECT 154.160 40.760 154.420 40.790 ;
        RECT 154.160 40.470 154.440 40.760 ;
        RECT 154.600 40.670 155.600 41.220 ;
        RECT 156.470 40.790 157.200 42.140 ;
        RECT 159.690 41.560 160.040 43.390 ;
        RECT 157.920 41.290 160.040 41.560 ;
        RECT 154.600 40.500 155.600 40.510 ;
        RECT 154.160 40.450 154.420 40.470 ;
        RECT 154.590 40.290 155.600 40.500 ;
        RECT 155.740 40.460 157.770 40.790 ;
        RECT 157.930 40.760 158.960 41.290 ;
        RECT 157.945 40.730 158.945 40.760 ;
        RECT 157.945 40.500 158.945 40.520 ;
        RECT 154.590 40.200 155.740 40.290 ;
        RECT 157.920 40.200 158.960 40.500 ;
        RECT 159.120 40.460 159.440 40.790 ;
        RECT 154.590 40.060 158.960 40.200 ;
        RECT 154.590 40.040 157.970 40.060 ;
        RECT 153.540 39.120 155.600 39.390 ;
        RECT 153.540 37.290 153.910 39.120 ;
        RECT 154.160 38.660 154.420 38.690 ;
        RECT 154.160 38.370 154.440 38.660 ;
        RECT 154.600 38.570 155.600 39.120 ;
        RECT 156.470 38.690 157.200 40.040 ;
        RECT 159.690 39.460 160.040 41.290 ;
        RECT 157.920 39.190 160.040 39.460 ;
        RECT 154.600 38.400 155.600 38.410 ;
        RECT 154.160 38.350 154.420 38.370 ;
        RECT 154.590 38.190 155.600 38.400 ;
        RECT 155.740 38.360 157.770 38.690 ;
        RECT 157.930 38.660 158.960 39.190 ;
        RECT 157.945 38.630 158.945 38.660 ;
        RECT 157.945 38.400 158.945 38.420 ;
        RECT 154.590 38.100 155.740 38.190 ;
        RECT 157.920 38.100 158.960 38.400 ;
        RECT 159.120 38.360 159.440 38.690 ;
        RECT 154.590 37.960 158.960 38.100 ;
        RECT 154.590 37.940 157.970 37.960 ;
        RECT 153.540 37.020 155.600 37.290 ;
        RECT 153.540 35.190 153.910 37.020 ;
        RECT 154.160 36.560 154.420 36.590 ;
        RECT 154.160 36.270 154.440 36.560 ;
        RECT 154.600 36.470 155.600 37.020 ;
        RECT 156.470 36.590 157.200 37.940 ;
        RECT 159.690 37.360 160.040 39.190 ;
        RECT 157.920 37.090 160.040 37.360 ;
        RECT 154.600 36.300 155.600 36.310 ;
        RECT 154.160 36.250 154.420 36.270 ;
        RECT 154.590 36.090 155.600 36.300 ;
        RECT 155.740 36.260 157.770 36.590 ;
        RECT 157.930 36.560 158.960 37.090 ;
        RECT 157.945 36.530 158.945 36.560 ;
        RECT 157.945 36.300 158.945 36.320 ;
        RECT 154.590 36.000 155.740 36.090 ;
        RECT 157.920 36.000 158.960 36.300 ;
        RECT 159.120 36.260 159.440 36.590 ;
        RECT 154.590 35.860 158.960 36.000 ;
        RECT 154.590 35.840 157.970 35.860 ;
        RECT 153.540 34.920 155.600 35.190 ;
        RECT 153.540 33.090 153.910 34.920 ;
        RECT 154.160 34.460 154.420 34.490 ;
        RECT 154.160 34.170 154.440 34.460 ;
        RECT 154.600 34.370 155.600 34.920 ;
        RECT 156.470 34.490 157.200 35.840 ;
        RECT 159.690 35.260 160.040 37.090 ;
        RECT 157.920 34.990 160.040 35.260 ;
        RECT 154.600 34.200 155.600 34.210 ;
        RECT 154.160 34.150 154.420 34.170 ;
        RECT 154.590 33.990 155.600 34.200 ;
        RECT 155.740 34.160 157.770 34.490 ;
        RECT 157.930 34.460 158.960 34.990 ;
        RECT 157.945 34.430 158.945 34.460 ;
        RECT 157.945 34.200 158.945 34.220 ;
        RECT 154.590 33.900 155.740 33.990 ;
        RECT 157.920 33.900 158.960 34.200 ;
        RECT 159.120 34.160 159.440 34.490 ;
        RECT 154.590 33.760 158.960 33.900 ;
        RECT 154.590 33.740 157.970 33.760 ;
        RECT 153.540 32.820 155.600 33.090 ;
        RECT 153.540 30.990 153.910 32.820 ;
        RECT 154.160 32.360 154.420 32.390 ;
        RECT 154.160 32.070 154.440 32.360 ;
        RECT 154.600 32.270 155.600 32.820 ;
        RECT 156.470 32.390 157.200 33.740 ;
        RECT 159.690 33.160 160.040 34.990 ;
        RECT 157.920 32.890 160.040 33.160 ;
        RECT 154.600 32.100 155.600 32.110 ;
        RECT 154.160 32.050 154.420 32.070 ;
        RECT 154.590 31.890 155.600 32.100 ;
        RECT 155.740 32.060 157.770 32.390 ;
        RECT 157.930 32.360 158.960 32.890 ;
        RECT 157.945 32.330 158.945 32.360 ;
        RECT 157.945 32.100 158.945 32.120 ;
        RECT 154.590 31.800 155.740 31.890 ;
        RECT 157.920 31.800 158.960 32.100 ;
        RECT 159.120 32.060 159.440 32.390 ;
        RECT 154.590 31.660 158.960 31.800 ;
        RECT 154.590 31.640 157.970 31.660 ;
        RECT 153.540 30.720 155.600 30.990 ;
        RECT 153.540 28.890 153.910 30.720 ;
        RECT 154.160 30.260 154.420 30.290 ;
        RECT 154.160 29.970 154.440 30.260 ;
        RECT 154.600 30.170 155.600 30.720 ;
        RECT 156.470 30.290 157.200 31.640 ;
        RECT 159.690 31.060 160.040 32.890 ;
        RECT 157.920 30.790 160.040 31.060 ;
        RECT 154.600 30.000 155.600 30.010 ;
        RECT 154.160 29.950 154.420 29.970 ;
        RECT 154.590 29.790 155.600 30.000 ;
        RECT 155.740 29.960 157.770 30.290 ;
        RECT 157.930 30.260 158.960 30.790 ;
        RECT 157.945 30.230 158.945 30.260 ;
        RECT 157.945 30.000 158.945 30.020 ;
        RECT 154.590 29.700 155.740 29.790 ;
        RECT 157.920 29.700 158.960 30.000 ;
        RECT 159.120 29.960 159.440 30.290 ;
        RECT 154.590 29.560 158.960 29.700 ;
        RECT 154.590 29.540 157.970 29.560 ;
        RECT 153.540 28.620 155.600 28.890 ;
        RECT 153.540 26.790 153.910 28.620 ;
        RECT 154.160 28.160 154.420 28.190 ;
        RECT 154.160 27.870 154.440 28.160 ;
        RECT 154.600 28.070 155.600 28.620 ;
        RECT 156.470 28.190 157.200 29.540 ;
        RECT 159.690 28.960 160.040 30.790 ;
        RECT 157.920 28.690 160.040 28.960 ;
        RECT 154.600 27.900 155.600 27.910 ;
        RECT 154.160 27.850 154.420 27.870 ;
        RECT 154.590 27.690 155.600 27.900 ;
        RECT 155.740 27.860 157.770 28.190 ;
        RECT 157.930 28.160 158.960 28.690 ;
        RECT 157.945 28.130 158.945 28.160 ;
        RECT 157.945 27.900 158.945 27.920 ;
        RECT 154.590 27.600 155.740 27.690 ;
        RECT 157.920 27.600 158.960 27.900 ;
        RECT 159.120 27.860 159.440 28.190 ;
        RECT 154.590 27.460 158.960 27.600 ;
        RECT 154.590 27.440 157.970 27.460 ;
        RECT 153.540 26.520 155.600 26.790 ;
        RECT 153.540 24.690 153.910 26.520 ;
        RECT 154.160 26.060 154.420 26.090 ;
        RECT 154.160 25.770 154.440 26.060 ;
        RECT 154.600 25.970 155.600 26.520 ;
        RECT 156.470 26.090 157.200 27.440 ;
        RECT 159.690 26.860 160.040 28.690 ;
        RECT 157.920 26.590 160.040 26.860 ;
        RECT 154.600 25.800 155.600 25.810 ;
        RECT 154.160 25.750 154.420 25.770 ;
        RECT 154.590 25.590 155.600 25.800 ;
        RECT 155.740 25.760 157.770 26.090 ;
        RECT 157.930 26.060 158.960 26.590 ;
        RECT 157.945 26.030 158.945 26.060 ;
        RECT 157.945 25.800 158.945 25.820 ;
        RECT 154.590 25.500 155.740 25.590 ;
        RECT 157.920 25.500 158.960 25.800 ;
        RECT 159.120 25.760 159.440 26.090 ;
        RECT 154.590 25.360 158.960 25.500 ;
        RECT 154.590 25.340 157.970 25.360 ;
        RECT 153.540 24.420 155.600 24.690 ;
        RECT 153.540 22.590 153.910 24.420 ;
        RECT 154.160 23.960 154.420 23.990 ;
        RECT 154.160 23.670 154.440 23.960 ;
        RECT 154.600 23.870 155.600 24.420 ;
        RECT 156.470 23.990 157.200 25.340 ;
        RECT 159.690 24.760 160.040 26.590 ;
        RECT 157.920 24.490 160.040 24.760 ;
        RECT 154.600 23.700 155.600 23.710 ;
        RECT 154.160 23.650 154.420 23.670 ;
        RECT 154.590 23.490 155.600 23.700 ;
        RECT 155.740 23.660 157.770 23.990 ;
        RECT 157.930 23.960 158.960 24.490 ;
        RECT 157.945 23.930 158.945 23.960 ;
        RECT 157.945 23.700 158.945 23.720 ;
        RECT 154.590 23.400 155.740 23.490 ;
        RECT 157.920 23.400 158.960 23.700 ;
        RECT 159.120 23.660 159.440 23.990 ;
        RECT 154.590 23.260 158.960 23.400 ;
        RECT 154.590 23.240 157.970 23.260 ;
        RECT 153.540 22.320 155.600 22.590 ;
        RECT 153.540 20.490 153.910 22.320 ;
        RECT 154.160 21.860 154.420 21.890 ;
        RECT 154.160 21.570 154.440 21.860 ;
        RECT 154.600 21.770 155.600 22.320 ;
        RECT 156.470 21.890 157.200 23.240 ;
        RECT 159.690 22.660 160.040 24.490 ;
        RECT 157.920 22.390 160.040 22.660 ;
        RECT 154.600 21.600 155.600 21.610 ;
        RECT 154.160 21.550 154.420 21.570 ;
        RECT 154.590 21.390 155.600 21.600 ;
        RECT 155.740 21.560 157.770 21.890 ;
        RECT 157.930 21.860 158.960 22.390 ;
        RECT 157.945 21.830 158.945 21.860 ;
        RECT 157.945 21.600 158.945 21.620 ;
        RECT 154.590 21.300 155.740 21.390 ;
        RECT 157.920 21.300 158.960 21.600 ;
        RECT 159.120 21.560 159.440 21.890 ;
        RECT 154.590 21.160 158.960 21.300 ;
        RECT 154.590 21.140 157.970 21.160 ;
        RECT 153.540 20.220 155.600 20.490 ;
        RECT 153.540 18.390 153.910 20.220 ;
        RECT 154.160 19.760 154.420 19.790 ;
        RECT 154.160 19.470 154.440 19.760 ;
        RECT 154.600 19.670 155.600 20.220 ;
        RECT 156.470 19.790 157.200 21.140 ;
        RECT 159.690 20.560 160.040 22.390 ;
        RECT 157.920 20.290 160.040 20.560 ;
        RECT 154.600 19.500 155.600 19.510 ;
        RECT 154.160 19.450 154.420 19.470 ;
        RECT 154.590 19.290 155.600 19.500 ;
        RECT 155.740 19.460 157.770 19.790 ;
        RECT 157.930 19.760 158.960 20.290 ;
        RECT 157.945 19.730 158.945 19.760 ;
        RECT 157.945 19.500 158.945 19.520 ;
        RECT 154.590 19.200 155.740 19.290 ;
        RECT 157.920 19.200 158.960 19.500 ;
        RECT 159.120 19.460 159.440 19.790 ;
        RECT 154.590 19.060 158.960 19.200 ;
        RECT 154.590 19.040 157.970 19.060 ;
        RECT 153.540 18.120 155.600 18.390 ;
        RECT 153.540 16.290 153.910 18.120 ;
        RECT 154.160 17.660 154.420 17.690 ;
        RECT 154.160 17.370 154.440 17.660 ;
        RECT 154.600 17.570 155.600 18.120 ;
        RECT 156.470 17.690 157.200 19.040 ;
        RECT 159.690 18.460 160.040 20.290 ;
        RECT 157.920 18.190 160.040 18.460 ;
        RECT 154.600 17.400 155.600 17.410 ;
        RECT 154.160 17.350 154.420 17.370 ;
        RECT 154.590 17.190 155.600 17.400 ;
        RECT 155.740 17.360 157.770 17.690 ;
        RECT 157.930 17.660 158.960 18.190 ;
        RECT 157.945 17.630 158.945 17.660 ;
        RECT 157.945 17.400 158.945 17.420 ;
        RECT 154.590 17.100 155.740 17.190 ;
        RECT 157.920 17.100 158.960 17.400 ;
        RECT 159.120 17.360 159.440 17.690 ;
        RECT 154.590 16.960 158.960 17.100 ;
        RECT 154.590 16.940 157.970 16.960 ;
        RECT 153.540 16.020 155.600 16.290 ;
        RECT 153.540 14.190 153.910 16.020 ;
        RECT 154.160 15.560 154.420 15.590 ;
        RECT 154.160 15.270 154.440 15.560 ;
        RECT 154.600 15.470 155.600 16.020 ;
        RECT 156.470 15.590 157.200 16.940 ;
        RECT 159.690 16.360 160.040 18.190 ;
        RECT 157.920 16.090 160.040 16.360 ;
        RECT 154.600 15.300 155.600 15.310 ;
        RECT 154.160 15.250 154.420 15.270 ;
        RECT 154.590 15.090 155.600 15.300 ;
        RECT 155.740 15.260 157.770 15.590 ;
        RECT 157.930 15.560 158.960 16.090 ;
        RECT 157.945 15.530 158.945 15.560 ;
        RECT 157.945 15.300 158.945 15.320 ;
        RECT 154.590 15.000 155.740 15.090 ;
        RECT 157.920 15.000 158.960 15.300 ;
        RECT 159.120 15.260 159.440 15.590 ;
        RECT 154.590 14.860 158.960 15.000 ;
        RECT 154.590 14.840 157.970 14.860 ;
        RECT 153.540 13.920 155.600 14.190 ;
        RECT 153.540 12.090 153.910 13.920 ;
        RECT 154.160 13.460 154.420 13.490 ;
        RECT 154.160 13.170 154.440 13.460 ;
        RECT 154.600 13.370 155.600 13.920 ;
        RECT 156.470 13.490 157.200 14.840 ;
        RECT 159.690 14.260 160.040 16.090 ;
        RECT 157.920 13.990 160.040 14.260 ;
        RECT 154.600 13.200 155.600 13.210 ;
        RECT 154.160 13.150 154.420 13.170 ;
        RECT 154.590 12.990 155.600 13.200 ;
        RECT 155.740 13.160 157.770 13.490 ;
        RECT 157.930 13.460 158.960 13.990 ;
        RECT 157.945 13.430 158.945 13.460 ;
        RECT 157.945 13.200 158.945 13.220 ;
        RECT 154.590 12.900 155.740 12.990 ;
        RECT 157.920 12.900 158.960 13.200 ;
        RECT 159.120 13.160 159.440 13.490 ;
        RECT 154.590 12.760 158.960 12.900 ;
        RECT 154.590 12.740 157.970 12.760 ;
        RECT 153.540 11.820 155.600 12.090 ;
        RECT 153.540 9.990 153.910 11.820 ;
        RECT 154.160 11.360 154.420 11.390 ;
        RECT 154.160 11.070 154.440 11.360 ;
        RECT 154.600 11.270 155.600 11.820 ;
        RECT 156.470 11.390 157.200 12.740 ;
        RECT 159.690 12.160 160.040 13.990 ;
        RECT 157.920 11.890 160.040 12.160 ;
        RECT 154.600 11.100 155.600 11.110 ;
        RECT 154.160 11.050 154.420 11.070 ;
        RECT 154.590 10.890 155.600 11.100 ;
        RECT 155.740 11.060 157.770 11.390 ;
        RECT 157.930 11.360 158.960 11.890 ;
        RECT 157.945 11.330 158.945 11.360 ;
        RECT 157.945 11.100 158.945 11.120 ;
        RECT 154.590 10.800 155.740 10.890 ;
        RECT 157.920 10.800 158.960 11.100 ;
        RECT 159.120 11.060 159.440 11.390 ;
        RECT 154.590 10.660 158.960 10.800 ;
        RECT 154.590 10.640 157.970 10.660 ;
        RECT 153.540 9.720 155.600 9.990 ;
        RECT 153.540 7.890 153.910 9.720 ;
        RECT 154.160 9.260 154.420 9.290 ;
        RECT 154.160 8.970 154.440 9.260 ;
        RECT 154.600 9.170 155.600 9.720 ;
        RECT 156.470 9.290 157.200 10.640 ;
        RECT 159.690 10.060 160.040 11.890 ;
        RECT 157.920 9.790 160.040 10.060 ;
        RECT 154.600 9.000 155.600 9.010 ;
        RECT 154.160 8.950 154.420 8.970 ;
        RECT 154.590 8.790 155.600 9.000 ;
        RECT 155.740 8.960 157.770 9.290 ;
        RECT 157.930 9.260 158.960 9.790 ;
        RECT 157.945 9.230 158.945 9.260 ;
        RECT 157.945 9.000 158.945 9.020 ;
        RECT 154.590 8.700 155.740 8.790 ;
        RECT 157.920 8.700 158.960 9.000 ;
        RECT 159.120 8.960 159.440 9.290 ;
        RECT 154.590 8.560 158.960 8.700 ;
        RECT 154.590 8.540 157.970 8.560 ;
        RECT 153.540 7.620 155.600 7.890 ;
        RECT 153.540 5.790 153.910 7.620 ;
        RECT 154.160 7.160 154.420 7.190 ;
        RECT 154.160 6.870 154.440 7.160 ;
        RECT 154.600 7.070 155.600 7.620 ;
        RECT 156.470 7.190 157.200 8.540 ;
        RECT 159.690 7.960 160.040 9.790 ;
        RECT 157.920 7.690 160.040 7.960 ;
        RECT 154.600 6.900 155.600 6.910 ;
        RECT 154.160 6.850 154.420 6.870 ;
        RECT 154.590 6.690 155.600 6.900 ;
        RECT 155.740 6.860 157.770 7.190 ;
        RECT 157.930 7.160 158.960 7.690 ;
        RECT 157.945 7.130 158.945 7.160 ;
        RECT 157.945 6.900 158.945 6.920 ;
        RECT 154.590 6.600 155.740 6.690 ;
        RECT 157.920 6.600 158.960 6.900 ;
        RECT 159.120 6.860 159.440 7.190 ;
        RECT 154.590 6.460 158.960 6.600 ;
        RECT 154.590 6.440 157.970 6.460 ;
        RECT 153.540 5.520 155.600 5.790 ;
        RECT 153.540 3.690 153.910 5.520 ;
        RECT 154.160 5.060 154.420 5.090 ;
        RECT 154.160 4.770 154.440 5.060 ;
        RECT 154.600 4.970 155.600 5.520 ;
        RECT 156.470 5.090 157.200 6.440 ;
        RECT 159.690 5.860 160.040 7.690 ;
        RECT 157.920 5.590 160.040 5.860 ;
        RECT 154.600 4.800 155.600 4.810 ;
        RECT 154.160 4.750 154.420 4.770 ;
        RECT 154.590 4.590 155.600 4.800 ;
        RECT 155.740 4.760 157.770 5.090 ;
        RECT 157.930 5.060 158.960 5.590 ;
        RECT 157.945 5.030 158.945 5.060 ;
        RECT 157.945 4.800 158.945 4.820 ;
        RECT 154.590 4.500 155.740 4.590 ;
        RECT 157.920 4.500 158.960 4.800 ;
        RECT 159.120 4.760 159.440 5.090 ;
        RECT 154.590 4.360 158.960 4.500 ;
        RECT 154.590 4.340 157.970 4.360 ;
        RECT 153.540 3.420 155.600 3.690 ;
        RECT 153.540 1.760 153.910 3.420 ;
        RECT 154.160 2.960 154.420 2.990 ;
        RECT 154.160 2.670 154.440 2.960 ;
        RECT 154.600 2.870 155.600 3.420 ;
        RECT 156.470 2.990 157.200 4.340 ;
        RECT 159.690 3.760 160.040 5.590 ;
        RECT 157.920 3.490 160.040 3.760 ;
        RECT 154.600 2.700 155.600 2.710 ;
        RECT 154.160 2.650 154.420 2.670 ;
        RECT 154.590 2.490 155.600 2.700 ;
        RECT 155.740 2.660 157.770 2.990 ;
        RECT 157.930 2.960 158.960 3.490 ;
        RECT 157.945 2.930 158.945 2.960 ;
        RECT 157.945 2.700 158.945 2.720 ;
        RECT 154.590 2.400 155.740 2.490 ;
        RECT 157.920 2.400 158.960 2.700 ;
        RECT 159.120 2.660 159.440 2.990 ;
        RECT 154.590 2.260 158.960 2.400 ;
        RECT 154.590 2.240 157.970 2.260 ;
        RECT 156.470 1.860 157.200 2.240 ;
        RECT 156.470 1.760 157.210 1.860 ;
        RECT 159.690 1.760 160.040 3.490 ;
        RECT 134.330 0.940 135.230 1.590 ;
        RECT 156.480 1.570 157.210 1.760 ;
        RECT 156.410 0.960 157.310 1.570 ;
      LAYER via ;
        RECT 14.170 212.190 19.560 214.510 ;
        RECT 131.300 211.930 131.930 212.680 ;
        RECT 134.540 210.540 135.070 211.610 ;
        RECT 153.230 212.100 154.170 212.580 ;
        RECT 134.470 1.880 135.100 2.290 ;
        RECT 156.550 210.730 157.080 211.680 ;
        RECT 156.540 1.890 157.100 2.320 ;
        RECT 134.430 1.070 135.160 1.470 ;
        RECT 156.510 1.070 157.220 1.460 ;
      LAYER met2 ;
        RECT 52.520 216.280 55.950 217.060 ;
        RECT 52.520 216.270 153.390 216.280 ;
        RECT 13.740 211.680 19.920 215.050 ;
        RECT 52.520 214.920 154.080 216.270 ;
        RECT 52.520 214.310 55.950 214.920 ;
        RECT 131.450 212.720 131.830 214.920 ;
        RECT 131.250 211.870 131.970 212.720 ;
        RECT 153.350 212.650 154.080 214.920 ;
        RECT 153.170 212.010 154.290 212.650 ;
        RECT 134.410 1.750 135.150 211.690 ;
        RECT 156.470 1.760 157.200 211.760 ;
        RECT 134.330 0.940 135.230 1.590 ;
        RECT 156.410 0.960 157.310 1.570 ;
      LAYER via2 ;
        RECT 14.170 212.190 19.560 214.510 ;
        RECT 52.840 214.800 55.520 216.700 ;
        RECT 134.430 1.070 135.160 1.470 ;
        RECT 156.510 1.070 157.220 1.460 ;
      LAYER met3 ;
        RECT 13.740 211.680 19.920 215.050 ;
        RECT 52.520 214.310 55.950 217.060 ;
        RECT 134.330 0.940 135.230 1.590 ;
        RECT 156.410 0.960 157.310 1.570 ;
      LAYER via3 ;
        RECT 14.170 212.190 19.560 214.510 ;
        RECT 52.840 214.800 55.520 216.700 ;
        RECT 134.430 1.070 135.160 1.470 ;
        RECT 156.510 1.070 157.220 1.460 ;
      LAYER met4 ;
        RECT 4.290 224.760 7.670 224.830 ;
        RECT 7.970 224.760 11.350 224.830 ;
        RECT 11.650 224.760 15.030 224.830 ;
        RECT 15.330 224.760 18.710 224.830 ;
        RECT 19.010 224.760 22.390 224.830 ;
        RECT 22.690 224.760 26.070 224.830 ;
        RECT 26.370 224.760 29.750 224.830 ;
        RECT 30.050 224.760 33.430 224.830 ;
        RECT 33.730 224.760 37.110 224.830 ;
        RECT 37.410 224.760 40.790 224.830 ;
        RECT 41.090 224.760 44.470 224.830 ;
        RECT 44.770 224.760 48.150 224.830 ;
        RECT 48.450 224.760 51.830 224.830 ;
        RECT 52.130 224.760 55.510 224.830 ;
        RECT 55.810 224.760 59.190 224.830 ;
        RECT 59.490 224.760 62.870 224.830 ;
        RECT 63.170 224.760 66.550 224.830 ;
        RECT 66.850 224.760 70.230 224.830 ;
        RECT 70.530 224.760 73.910 224.830 ;
        RECT 74.210 224.760 77.590 224.830 ;
        RECT 77.890 224.760 81.270 224.830 ;
        RECT 81.570 224.760 84.950 224.830 ;
        RECT 85.250 224.760 88.630 224.830 ;
        RECT 88.930 224.760 88.940 224.830 ;
        RECT 3.990 222.480 88.940 224.760 ;
        RECT 49.000 220.760 50.500 222.480 ;
        RECT 52.520 216.290 55.950 217.060 ;
        RECT 13.740 213.960 19.920 215.050 ;
        RECT 50.500 214.920 55.950 216.290 ;
        RECT 52.520 214.310 55.950 214.920 ;
        RECT 2.500 212.920 19.920 213.960 ;
        RECT 13.740 211.680 19.920 212.920 ;
        RECT 134.330 1.000 135.230 1.590 ;
        RECT 156.410 1.000 157.310 1.570 ;
  END
END tt_um_devin
END LIBRARY

